// $Header: $
///////////////////////////////////////////////////////
//  Copyright (c) 2011 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /     Vendor      : Xilinx 
// \  \    \/      Version     :  13.1
//  \  \           Description : 
//  /  /                      
// /__/   /\       Filename    : PCIE_3_0.uniprim.v
// \  \  /  \ 
//  \__\/\__ \                    
//                                 
//  Generated by :	/home/chen/xfoundry/HEAD/env/Databases/CAEInterfaces/LibraryWriters/bin/ltw.pl
//  Revision:		1.0
//  01/18/13 - 695630 - added drp monitor
///////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

`celldefine

module PCIE_3_0 (
  CFGCURRENTSPEED,
  CFGDPASUBSTATECHANGE,
  CFGERRCOROUT,
  CFGERRFATALOUT,
  CFGERRNONFATALOUT,
  CFGEXTFUNCTIONNUMBER,
  CFGEXTREADRECEIVED,
  CFGEXTREGISTERNUMBER,
  CFGEXTWRITEBYTEENABLE,
  CFGEXTWRITEDATA,
  CFGEXTWRITERECEIVED,
  CFGFCCPLD,
  CFGFCCPLH,
  CFGFCNPD,
  CFGFCNPH,
  CFGFCPD,
  CFGFCPH,
  CFGFLRINPROCESS,
  CFGFUNCTIONPOWERSTATE,
  CFGFUNCTIONSTATUS,
  CFGHOTRESETOUT,
  CFGINPUTUPDATEDONE,
  CFGINTERRUPTAOUTPUT,
  CFGINTERRUPTBOUTPUT,
  CFGINTERRUPTCOUTPUT,
  CFGINTERRUPTDOUTPUT,
  CFGINTERRUPTMSIDATA,
  CFGINTERRUPTMSIENABLE,
  CFGINTERRUPTMSIFAIL,
  CFGINTERRUPTMSIMASKUPDATE,
  CFGINTERRUPTMSIMMENABLE,
  CFGINTERRUPTMSISENT,
  CFGINTERRUPTMSIVFENABLE,
  CFGINTERRUPTMSIXENABLE,
  CFGINTERRUPTMSIXFAIL,
  CFGINTERRUPTMSIXMASK,
  CFGINTERRUPTMSIXSENT,
  CFGINTERRUPTMSIXVFENABLE,
  CFGINTERRUPTMSIXVFMASK,
  CFGINTERRUPTSENT,
  CFGLINKPOWERSTATE,
  CFGLOCALERROR,
  CFGLTRENABLE,
  CFGLTSSMSTATE,
  CFGMAXPAYLOAD,
  CFGMAXREADREQ,
  CFGMCUPDATEDONE,
  CFGMGMTREADDATA,
  CFGMGMTREADWRITEDONE,
  CFGMSGRECEIVED,
  CFGMSGRECEIVEDDATA,
  CFGMSGRECEIVEDTYPE,
  CFGMSGTRANSMITDONE,
  CFGNEGOTIATEDWIDTH,
  CFGOBFFENABLE,
  CFGPERFUNCSTATUSDATA,
  CFGPERFUNCTIONUPDATEDONE,
  CFGPHYLINKDOWN,
  CFGPHYLINKSTATUS,
  CFGPLSTATUSCHANGE,
  CFGPOWERSTATECHANGEINTERRUPT,
  CFGRCBSTATUS,
  CFGTPHFUNCTIONNUM,
  CFGTPHREQUESTERENABLE,
  CFGTPHSTMODE,
  CFGTPHSTTADDRESS,
  CFGTPHSTTREADENABLE,
  CFGTPHSTTWRITEBYTEVALID,
  CFGTPHSTTWRITEDATA,
  CFGTPHSTTWRITEENABLE,
  CFGVFFLRINPROCESS,
  CFGVFPOWERSTATE,
  CFGVFSTATUS,
  CFGVFTPHREQUESTERENABLE,
  CFGVFTPHSTMODE,
  DBGDATAOUT,
  DRPDO,
  DRPRDY,
  MAXISCQTDATA,
  MAXISCQTKEEP,
  MAXISCQTLAST,
  MAXISCQTUSER,
  MAXISCQTVALID,
  MAXISRCTDATA,
  MAXISRCTKEEP,
  MAXISRCTLAST,
  MAXISRCTUSER,
  MAXISRCTVALID,
  MICOMPLETIONRAMREADADDRESSAL,
  MICOMPLETIONRAMREADADDRESSAU,
  MICOMPLETIONRAMREADADDRESSBL,
  MICOMPLETIONRAMREADADDRESSBU,
  MICOMPLETIONRAMREADENABLEL,
  MICOMPLETIONRAMREADENABLEU,
  MICOMPLETIONRAMWRITEADDRESSAL,
  MICOMPLETIONRAMWRITEADDRESSAU,
  MICOMPLETIONRAMWRITEADDRESSBL,
  MICOMPLETIONRAMWRITEADDRESSBU,
  MICOMPLETIONRAMWRITEDATAL,
  MICOMPLETIONRAMWRITEDATAU,
  MICOMPLETIONRAMWRITEENABLEL,
  MICOMPLETIONRAMWRITEENABLEU,
  MIREPLAYRAMADDRESS,
  MIREPLAYRAMREADENABLE,
  MIREPLAYRAMWRITEDATA,
  MIREPLAYRAMWRITEENABLE,
  MIREQUESTRAMREADADDRESSA,
  MIREQUESTRAMREADADDRESSB,
  MIREQUESTRAMREADENABLE,
  MIREQUESTRAMWRITEADDRESSA,
  MIREQUESTRAMWRITEADDRESSB,
  MIREQUESTRAMWRITEDATA,
  MIREQUESTRAMWRITEENABLE,
  PCIECQNPREQCOUNT,
  PCIERQSEQNUM,
  PCIERQSEQNUMVLD,
  PCIERQTAG,
  PCIERQTAGAV,
  PCIERQTAGVLD,
  PCIETFCNPDAV,
  PCIETFCNPHAV,
  PIPERX0EQCONTROL,
  PIPERX0EQLPLFFS,
  PIPERX0EQLPTXPRESET,
  PIPERX0EQPRESET,
  PIPERX0POLARITY,
  PIPERX1EQCONTROL,
  PIPERX1EQLPLFFS,
  PIPERX1EQLPTXPRESET,
  PIPERX1EQPRESET,
  PIPERX1POLARITY,
  PIPERX2EQCONTROL,
  PIPERX2EQLPLFFS,
  PIPERX2EQLPTXPRESET,
  PIPERX2EQPRESET,
  PIPERX2POLARITY,
  PIPERX3EQCONTROL,
  PIPERX3EQLPLFFS,
  PIPERX3EQLPTXPRESET,
  PIPERX3EQPRESET,
  PIPERX3POLARITY,
  PIPERX4EQCONTROL,
  PIPERX4EQLPLFFS,
  PIPERX4EQLPTXPRESET,
  PIPERX4EQPRESET,
  PIPERX4POLARITY,
  PIPERX5EQCONTROL,
  PIPERX5EQLPLFFS,
  PIPERX5EQLPTXPRESET,
  PIPERX5EQPRESET,
  PIPERX5POLARITY,
  PIPERX6EQCONTROL,
  PIPERX6EQLPLFFS,
  PIPERX6EQLPTXPRESET,
  PIPERX6EQPRESET,
  PIPERX6POLARITY,
  PIPERX7EQCONTROL,
  PIPERX7EQLPLFFS,
  PIPERX7EQLPTXPRESET,
  PIPERX7EQPRESET,
  PIPERX7POLARITY,
  PIPETX0CHARISK,
  PIPETX0COMPLIANCE,
  PIPETX0DATA,
  PIPETX0DATAVALID,
  PIPETX0ELECIDLE,
  PIPETX0EQCONTROL,
  PIPETX0EQDEEMPH,
  PIPETX0EQPRESET,
  PIPETX0POWERDOWN,
  PIPETX0STARTBLOCK,
  PIPETX0SYNCHEADER,
  PIPETX1CHARISK,
  PIPETX1COMPLIANCE,
  PIPETX1DATA,
  PIPETX1DATAVALID,
  PIPETX1ELECIDLE,
  PIPETX1EQCONTROL,
  PIPETX1EQDEEMPH,
  PIPETX1EQPRESET,
  PIPETX1POWERDOWN,
  PIPETX1STARTBLOCK,
  PIPETX1SYNCHEADER,
  PIPETX2CHARISK,
  PIPETX2COMPLIANCE,
  PIPETX2DATA,
  PIPETX2DATAVALID,
  PIPETX2ELECIDLE,
  PIPETX2EQCONTROL,
  PIPETX2EQDEEMPH,
  PIPETX2EQPRESET,
  PIPETX2POWERDOWN,
  PIPETX2STARTBLOCK,
  PIPETX2SYNCHEADER,
  PIPETX3CHARISK,
  PIPETX3COMPLIANCE,
  PIPETX3DATA,
  PIPETX3DATAVALID,
  PIPETX3ELECIDLE,
  PIPETX3EQCONTROL,
  PIPETX3EQDEEMPH,
  PIPETX3EQPRESET,
  PIPETX3POWERDOWN,
  PIPETX3STARTBLOCK,
  PIPETX3SYNCHEADER,
  PIPETX4CHARISK,
  PIPETX4COMPLIANCE,
  PIPETX4DATA,
  PIPETX4DATAVALID,
  PIPETX4ELECIDLE,
  PIPETX4EQCONTROL,
  PIPETX4EQDEEMPH,
  PIPETX4EQPRESET,
  PIPETX4POWERDOWN,
  PIPETX4STARTBLOCK,
  PIPETX4SYNCHEADER,
  PIPETX5CHARISK,
  PIPETX5COMPLIANCE,
  PIPETX5DATA,
  PIPETX5DATAVALID,
  PIPETX5ELECIDLE,
  PIPETX5EQCONTROL,
  PIPETX5EQDEEMPH,
  PIPETX5EQPRESET,
  PIPETX5POWERDOWN,
  PIPETX5STARTBLOCK,
  PIPETX5SYNCHEADER,
  PIPETX6CHARISK,
  PIPETX6COMPLIANCE,
  PIPETX6DATA,
  PIPETX6DATAVALID,
  PIPETX6ELECIDLE,
  PIPETX6EQCONTROL,
  PIPETX6EQDEEMPH,
  PIPETX6EQPRESET,
  PIPETX6POWERDOWN,
  PIPETX6STARTBLOCK,
  PIPETX6SYNCHEADER,
  PIPETX7CHARISK,
  PIPETX7COMPLIANCE,
  PIPETX7DATA,
  PIPETX7DATAVALID,
  PIPETX7ELECIDLE,
  PIPETX7EQCONTROL,
  PIPETX7EQDEEMPH,
  PIPETX7EQPRESET,
  PIPETX7POWERDOWN,
  PIPETX7STARTBLOCK,
  PIPETX7SYNCHEADER,
  PIPETXDEEMPH,
  PIPETXMARGIN,
  PIPETXRATE,
  PIPETXRCVRDET,
  PIPETXRESET,
  PIPETXSWING,
  PLEQINPROGRESS,
  PLEQPHASE,
  PLGEN3PCSRXSLIDE,
  SAXISCCTREADY,
  SAXISRQTREADY,

  CFGCONFIGSPACEENABLE,
  CFGDEVID,
  CFGDSBUSNUMBER,
  CFGDSDEVICENUMBER,
  CFGDSFUNCTIONNUMBER,
  CFGDSN,
  CFGDSPORTNUMBER,
  CFGERRCORIN,
  CFGERRUNCORIN,
  CFGEXTREADDATA,
  CFGEXTREADDATAVALID,
  CFGFCSEL,
  CFGFLRDONE,
  CFGHOTRESETIN,
  CFGINPUTUPDATEREQUEST,
  CFGINTERRUPTINT,
  CFGINTERRUPTMSIATTR,
  CFGINTERRUPTMSIFUNCTIONNUMBER,
  CFGINTERRUPTMSIINT,
  CFGINTERRUPTMSIPENDINGSTATUS,
  CFGINTERRUPTMSISELECT,
  CFGINTERRUPTMSITPHPRESENT,
  CFGINTERRUPTMSITPHSTTAG,
  CFGINTERRUPTMSITPHTYPE,
  CFGINTERRUPTMSIXADDRESS,
  CFGINTERRUPTMSIXDATA,
  CFGINTERRUPTMSIXINT,
  CFGINTERRUPTPENDING,
  CFGLINKTRAININGENABLE,
  CFGMCUPDATEREQUEST,
  CFGMGMTADDR,
  CFGMGMTBYTEENABLE,
  CFGMGMTREAD,
  CFGMGMTTYPE1CFGREGACCESS,
  CFGMGMTWRITE,
  CFGMGMTWRITEDATA,
  CFGMSGTRANSMIT,
  CFGMSGTRANSMITDATA,
  CFGMSGTRANSMITTYPE,
  CFGPERFUNCSTATUSCONTROL,
  CFGPERFUNCTIONNUMBER,
  CFGPERFUNCTIONOUTPUTREQUEST,
  CFGPOWERSTATECHANGEACK,
  CFGREQPMTRANSITIONL23READY,
  CFGREVID,
  CFGSUBSYSID,
  CFGSUBSYSVENDID,
  CFGTPHSTTREADDATA,
  CFGTPHSTTREADDATAVALID,
  CFGVENDID,
  CFGVFFLRDONE,
  CORECLK,
  CORECLKMICOMPLETIONRAML,
  CORECLKMICOMPLETIONRAMU,
  CORECLKMIREPLAYRAM,
  CORECLKMIREQUESTRAM,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  MAXISCQTREADY,
  MAXISRCTREADY,
  MGMTRESETN,
  MGMTSTICKYRESETN,
  MICOMPLETIONRAMREADDATA,
  MIREPLAYRAMREADDATA,
  MIREQUESTRAMREADDATA,
  PCIECQNPREQ,
  PIPECLK,
  PIPEEQFS,
  PIPEEQLF,
  PIPERESETN,
  PIPERX0CHARISK,
  PIPERX0DATA,
  PIPERX0DATAVALID,
  PIPERX0ELECIDLE,
  PIPERX0EQDONE,
  PIPERX0EQLPADAPTDONE,
  PIPERX0EQLPLFFSSEL,
  PIPERX0EQLPNEWTXCOEFFORPRESET,
  PIPERX0PHYSTATUS,
  PIPERX0STARTBLOCK,
  PIPERX0STATUS,
  PIPERX0SYNCHEADER,
  PIPERX0VALID,
  PIPERX1CHARISK,
  PIPERX1DATA,
  PIPERX1DATAVALID,
  PIPERX1ELECIDLE,
  PIPERX1EQDONE,
  PIPERX1EQLPADAPTDONE,
  PIPERX1EQLPLFFSSEL,
  PIPERX1EQLPNEWTXCOEFFORPRESET,
  PIPERX1PHYSTATUS,
  PIPERX1STARTBLOCK,
  PIPERX1STATUS,
  PIPERX1SYNCHEADER,
  PIPERX1VALID,
  PIPERX2CHARISK,
  PIPERX2DATA,
  PIPERX2DATAVALID,
  PIPERX2ELECIDLE,
  PIPERX2EQDONE,
  PIPERX2EQLPADAPTDONE,
  PIPERX2EQLPLFFSSEL,
  PIPERX2EQLPNEWTXCOEFFORPRESET,
  PIPERX2PHYSTATUS,
  PIPERX2STARTBLOCK,
  PIPERX2STATUS,
  PIPERX2SYNCHEADER,
  PIPERX2VALID,
  PIPERX3CHARISK,
  PIPERX3DATA,
  PIPERX3DATAVALID,
  PIPERX3ELECIDLE,
  PIPERX3EQDONE,
  PIPERX3EQLPADAPTDONE,
  PIPERX3EQLPLFFSSEL,
  PIPERX3EQLPNEWTXCOEFFORPRESET,
  PIPERX3PHYSTATUS,
  PIPERX3STARTBLOCK,
  PIPERX3STATUS,
  PIPERX3SYNCHEADER,
  PIPERX3VALID,
  PIPERX4CHARISK,
  PIPERX4DATA,
  PIPERX4DATAVALID,
  PIPERX4ELECIDLE,
  PIPERX4EQDONE,
  PIPERX4EQLPADAPTDONE,
  PIPERX4EQLPLFFSSEL,
  PIPERX4EQLPNEWTXCOEFFORPRESET,
  PIPERX4PHYSTATUS,
  PIPERX4STARTBLOCK,
  PIPERX4STATUS,
  PIPERX4SYNCHEADER,
  PIPERX4VALID,
  PIPERX5CHARISK,
  PIPERX5DATA,
  PIPERX5DATAVALID,
  PIPERX5ELECIDLE,
  PIPERX5EQDONE,
  PIPERX5EQLPADAPTDONE,
  PIPERX5EQLPLFFSSEL,
  PIPERX5EQLPNEWTXCOEFFORPRESET,
  PIPERX5PHYSTATUS,
  PIPERX5STARTBLOCK,
  PIPERX5STATUS,
  PIPERX5SYNCHEADER,
  PIPERX5VALID,
  PIPERX6CHARISK,
  PIPERX6DATA,
  PIPERX6DATAVALID,
  PIPERX6ELECIDLE,
  PIPERX6EQDONE,
  PIPERX6EQLPADAPTDONE,
  PIPERX6EQLPLFFSSEL,
  PIPERX6EQLPNEWTXCOEFFORPRESET,
  PIPERX6PHYSTATUS,
  PIPERX6STARTBLOCK,
  PIPERX6STATUS,
  PIPERX6SYNCHEADER,
  PIPERX6VALID,
  PIPERX7CHARISK,
  PIPERX7DATA,
  PIPERX7DATAVALID,
  PIPERX7ELECIDLE,
  PIPERX7EQDONE,
  PIPERX7EQLPADAPTDONE,
  PIPERX7EQLPLFFSSEL,
  PIPERX7EQLPNEWTXCOEFFORPRESET,
  PIPERX7PHYSTATUS,
  PIPERX7STARTBLOCK,
  PIPERX7STATUS,
  PIPERX7SYNCHEADER,
  PIPERX7VALID,
  PIPETX0EQCOEFF,
  PIPETX0EQDONE,
  PIPETX1EQCOEFF,
  PIPETX1EQDONE,
  PIPETX2EQCOEFF,
  PIPETX2EQDONE,
  PIPETX3EQCOEFF,
  PIPETX3EQDONE,
  PIPETX4EQCOEFF,
  PIPETX4EQDONE,
  PIPETX5EQCOEFF,
  PIPETX5EQDONE,
  PIPETX6EQCOEFF,
  PIPETX6EQDONE,
  PIPETX7EQCOEFF,
  PIPETX7EQDONE,
  PLDISABLESCRAMBLER,
  PLEQRESETEIEOSCOUNT,
  PLGEN3PCSDISABLE,
  PLGEN3PCSRXSYNCDONE,
  RECCLK,
  RESETN,
  SAXISCCTDATA,
  SAXISCCTKEEP,
  SAXISCCTLAST,
  SAXISCCTUSER,
  SAXISCCTVALID,
  SAXISRQTDATA,
  SAXISRQTKEEP,
  SAXISRQTLAST,
  SAXISRQTUSER,
  SAXISRQTVALID,
  USERCLK
);

  `ifdef XIL_TIMING //Simprim 
  parameter LOC = "UNPLACED";
  `endif
  parameter ARI_CAP_ENABLE = "FALSE";
  parameter AXISTEN_IF_CC_ALIGNMENT_MODE = "FALSE";
  parameter AXISTEN_IF_CC_PARITY_CHK = "TRUE";
  parameter AXISTEN_IF_CQ_ALIGNMENT_MODE = "FALSE";
  parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
  parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
  parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
  parameter AXISTEN_IF_RC_ALIGNMENT_MODE = "FALSE";
  parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
  parameter AXISTEN_IF_RQ_ALIGNMENT_MODE = "FALSE";
  parameter AXISTEN_IF_RQ_PARITY_CHK = "TRUE";
  parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
  parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
  parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
  parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
  parameter [1:0] GEN3_PCS_AUTO_REALIGN = 2'h1;
  parameter GEN3_PCS_RX_ELECIDLE_INTERNAL = "TRUE";
  parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
  parameter LL_ACK_TIMEOUT_EN = "FALSE";
  parameter integer LL_ACK_TIMEOUT_FUNC = 0;
  parameter [15:0] LL_CPL_FC_UPDATE_TIMER = 16'h0000;
  parameter LL_CPL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
  parameter [15:0] LL_FC_UPDATE_TIMER = 16'h0000;
  parameter LL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
  parameter [15:0] LL_NP_FC_UPDATE_TIMER = 16'h0000;
  parameter LL_NP_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
  parameter [15:0] LL_P_FC_UPDATE_TIMER = 16'h0000;
  parameter LL_P_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
  parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
  parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
  parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
  parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h0FA;
  parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
  parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
  parameter PF0_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
  parameter PF0_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
  parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
  parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
  parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
  parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
  parameter [4:0] PF0_BAR0_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
  parameter [4:0] PF0_BAR1_APERTURE_SIZE = 5'h00;
  parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
  parameter [4:0] PF0_BAR2_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
  parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
  parameter [4:0] PF0_BAR4_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
  parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
  parameter [7:0] PF0_BIST_REGISTER = 8'h00;
  parameter [7:0] PF0_CAPABILITY_POINTER = 8'h50;
  parameter [23:0] PF0_CLASS_CODE = 24'h000000;
  parameter [15:0] PF0_DEVICE_ID = 16'h0000;
  parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
  parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
  parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
  parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
  parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
  parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
  parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
  parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
  parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
  parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
  parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
  parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
  parameter [11:0] PF0_DPA_CAP_NEXTPTR = 12'h000;
  parameter [4:0] PF0_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
  parameter PF0_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
  parameter [3:0] PF0_DPA_CAP_VER = 4'h1;
  parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
  parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
  parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
  parameter [7:0] PF0_INTERRUPT_LINE = 8'h00;
  parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
  parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
  parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
  parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
  parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
  parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
  parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
  parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
  parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
  parameter [11:0] PF0_PB_CAP_NEXTPTR = 12'h000;
  parameter PF0_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
  parameter [3:0] PF0_PB_CAP_VER = 4'h1;
  parameter [7:0] PF0_PM_CAP_ID = 8'h01;
  parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
  parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
  parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
  parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
  parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
  parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
  parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
  parameter PF0_RBAR_CAP_ENABLE = "FALSE";
  parameter [2:0] PF0_RBAR_CAP_INDEX0 = 3'h0;
  parameter [2:0] PF0_RBAR_CAP_INDEX1 = 3'h0;
  parameter [2:0] PF0_RBAR_CAP_INDEX2 = 3'h0;
  parameter [11:0] PF0_RBAR_CAP_NEXTPTR = 12'h000;
  parameter [19:0] PF0_RBAR_CAP_SIZE0 = 20'h00000;
  parameter [19:0] PF0_RBAR_CAP_SIZE1 = 20'h00000;
  parameter [19:0] PF0_RBAR_CAP_SIZE2 = 20'h00000;
  parameter [3:0] PF0_RBAR_CAP_VER = 4'h1;
  parameter [2:0] PF0_RBAR_NUM = 3'h1;
  parameter [7:0] PF0_REVISION_ID = 8'h00;
  parameter [4:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
  parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
  parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
  parameter [4:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
  parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
  parameter [4:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
  parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
  parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
  parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
  parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
  parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
  parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
  parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
  parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
  parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
  parameter [15:0] PF0_SUBSYSTEM_ID = 16'h0000;
  parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter PF0_TPHR_CAP_ENABLE = "FALSE";
  parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
  parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
  parameter [3:0] PF0_VC_CAP_VER = 4'h1;
  parameter PF1_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
  parameter PF1_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
  parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
  parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
  parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
  parameter [4:0] PF1_BAR0_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
  parameter [4:0] PF1_BAR1_APERTURE_SIZE = 5'h00;
  parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
  parameter [4:0] PF1_BAR2_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
  parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
  parameter [4:0] PF1_BAR4_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
  parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
  parameter [7:0] PF1_BIST_REGISTER = 8'h00;
  parameter [7:0] PF1_CAPABILITY_POINTER = 8'h50;
  parameter [23:0] PF1_CLASS_CODE = 24'h000000;
  parameter [15:0] PF1_DEVICE_ID = 16'h0000;
  parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
  parameter [11:0] PF1_DPA_CAP_NEXTPTR = 12'h000;
  parameter [4:0] PF1_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
  parameter PF1_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
  parameter [3:0] PF1_DPA_CAP_VER = 4'h1;
  parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
  parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
  parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
  parameter [7:0] PF1_INTERRUPT_LINE = 8'h00;
  parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
  parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
  parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
  parameter [11:0] PF1_PB_CAP_NEXTPTR = 12'h000;
  parameter PF1_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
  parameter [3:0] PF1_PB_CAP_VER = 4'h1;
  parameter [7:0] PF1_PM_CAP_ID = 8'h01;
  parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] PF1_PM_CAP_VER_ID = 3'h3;
  parameter PF1_RBAR_CAP_ENABLE = "FALSE";
  parameter [2:0] PF1_RBAR_CAP_INDEX0 = 3'h0;
  parameter [2:0] PF1_RBAR_CAP_INDEX1 = 3'h0;
  parameter [2:0] PF1_RBAR_CAP_INDEX2 = 3'h0;
  parameter [11:0] PF1_RBAR_CAP_NEXTPTR = 12'h000;
  parameter [19:0] PF1_RBAR_CAP_SIZE0 = 20'h00000;
  parameter [19:0] PF1_RBAR_CAP_SIZE1 = 20'h00000;
  parameter [19:0] PF1_RBAR_CAP_SIZE2 = 20'h00000;
  parameter [3:0] PF1_RBAR_CAP_VER = 4'h1;
  parameter [2:0] PF1_RBAR_NUM = 3'h1;
  parameter [7:0] PF1_REVISION_ID = 8'h00;
  parameter [4:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
  parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
  parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
  parameter [4:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
  parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
  parameter [4:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
  parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
  parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
  parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
  parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
  parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
  parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
  parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
  parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
  parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
  parameter [15:0] PF1_SUBSYSTEM_ID = 16'h0000;
  parameter PF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter PF1_TPHR_CAP_ENABLE = "FALSE";
  parameter PF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] PF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] PF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] PF1_TPHR_CAP_VER = 4'h1;
  parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
  parameter PL_DISABLE_GEN3_DC_BALANCE = "FALSE";
  parameter PL_DISABLE_SCRAMBLING = "FALSE";
  parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
  parameter PL_EQ_ADAPT_DISABLE_COEFF_CHECK = "FALSE";
  parameter PL_EQ_ADAPT_DISABLE_PRESET_CHECK = "FALSE";
  parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
  parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
  parameter PL_EQ_BYPASS_PHASE23 = "FALSE";
  parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
  parameter [15:0] PL_LANE0_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE1_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE2_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE3_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE4_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE5_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE6_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE7_EQ_CONTROL = 16'h3F00;
  parameter [2:0] PL_LINK_CAP_MAX_LINK_SPEED = 3'h4;
  parameter [3:0] PL_LINK_CAP_MAX_LINK_WIDTH = 4'h8;
  parameter integer PL_N_FTS_COMCLK_GEN1 = 255;
  parameter integer PL_N_FTS_COMCLK_GEN2 = 255;
  parameter integer PL_N_FTS_COMCLK_GEN3 = 255;
  parameter integer PL_N_FTS_GEN1 = 255;
  parameter integer PL_N_FTS_GEN2 = 255;
  parameter integer PL_N_FTS_GEN3 = 255;
  parameter PL_SIM_FAST_LINK_TRAINING = "FALSE";
  parameter PL_UPSTREAM_FACING = "TRUE";
  parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h05DC;
  parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h00000;
  parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
  parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000000;
  parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h186A0;
  parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0064;
  parameter SIM_VERSION = "1.0";
  parameter integer SPARE_BIT0 = 0;
  parameter integer SPARE_BIT1 = 0;
  parameter integer SPARE_BIT2 = 0;
  parameter integer SPARE_BIT3 = 0;
  parameter integer SPARE_BIT4 = 0;
  parameter integer SPARE_BIT5 = 0;
  parameter integer SPARE_BIT6 = 0;
  parameter integer SPARE_BIT7 = 0;
  parameter integer SPARE_BIT8 = 0;
  parameter [7:0] SPARE_BYTE0 = 8'h00;
  parameter [7:0] SPARE_BYTE1 = 8'h00;
  parameter [7:0] SPARE_BYTE2 = 8'h00;
  parameter [7:0] SPARE_BYTE3 = 8'h00;
  parameter [31:0] SPARE_WORD0 = 32'h00000000;
  parameter [31:0] SPARE_WORD1 = 32'h00000000;
  parameter [31:0] SPARE_WORD2 = 32'h00000000;
  parameter [31:0] SPARE_WORD3 = 32'h00000000;
  parameter SRIOV_CAP_ENABLE = "FALSE";
  parameter [23:0] TL_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
  parameter [27:0] TL_COMPL_TIMEOUT_REG1 = 28'h0000000;
  parameter [11:0] TL_CREDITS_CD = 12'h3E0;
  parameter [7:0] TL_CREDITS_CH = 8'h20;
  parameter [11:0] TL_CREDITS_NPD = 12'h028;
  parameter [7:0] TL_CREDITS_NPH = 8'h20;
  parameter [11:0] TL_CREDITS_PD = 12'h198;
  parameter [7:0] TL_CREDITS_PH = 8'h20;
  parameter TL_ENABLE_MESSAGE_RID_CHECK_ENABLE = "TRUE";
  parameter TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
  parameter TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
  parameter TL_LEGACY_MODE_ENABLE = "FALSE";
  parameter TL_PF_ENABLE_REG = "FALSE";
  parameter TL_TAG_MGMT_ENABLE = "TRUE";
  parameter [11:0] VF0_ARI_CAP_NEXTPTR = 12'h000;
  parameter [7:0] VF0_CAPABILITY_POINTER = 8'h50;
  parameter integer VF0_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF0_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF0_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF0_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF0_PM_CAP_ID = 8'h01;
  parameter [7:0] VF0_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF0_PM_CAP_VER_ID = 3'h3;
  parameter VF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF0_TPHR_CAP_ENABLE = "FALSE";
  parameter VF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF0_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF0_TPHR_CAP_VER = 4'h1;
  parameter [11:0] VF1_ARI_CAP_NEXTPTR = 12'h000;
  parameter integer VF1_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF1_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF1_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF1_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF1_PM_CAP_ID = 8'h01;
  parameter [7:0] VF1_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF1_PM_CAP_VER_ID = 3'h3;
  parameter VF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF1_TPHR_CAP_ENABLE = "FALSE";
  parameter VF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF1_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF1_TPHR_CAP_VER = 4'h1;
  parameter [11:0] VF2_ARI_CAP_NEXTPTR = 12'h000;
  parameter integer VF2_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF2_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF2_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF2_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF2_PM_CAP_ID = 8'h01;
  parameter [7:0] VF2_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF2_PM_CAP_VER_ID = 3'h3;
  parameter VF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF2_TPHR_CAP_ENABLE = "FALSE";
  parameter VF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF2_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF2_TPHR_CAP_VER = 4'h1;
  parameter [11:0] VF3_ARI_CAP_NEXTPTR = 12'h000;
  parameter integer VF3_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF3_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF3_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF3_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF3_PM_CAP_ID = 8'h01;
  parameter [7:0] VF3_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF3_PM_CAP_VER_ID = 3'h3;
  parameter VF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF3_TPHR_CAP_ENABLE = "FALSE";
  parameter VF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF3_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF3_TPHR_CAP_VER = 4'h1;
  parameter [11:0] VF4_ARI_CAP_NEXTPTR = 12'h000;
  parameter integer VF4_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF4_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF4_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF4_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF4_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF4_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF4_PM_CAP_ID = 8'h01;
  parameter [7:0] VF4_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF4_PM_CAP_VER_ID = 3'h3;
  parameter VF4_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF4_TPHR_CAP_ENABLE = "FALSE";
  parameter VF4_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF4_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF4_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF4_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF4_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF4_TPHR_CAP_VER = 4'h1;
  parameter [11:0] VF5_ARI_CAP_NEXTPTR = 12'h000;
  parameter integer VF5_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF5_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF5_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF5_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF5_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF5_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF5_PM_CAP_ID = 8'h01;
  parameter [7:0] VF5_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF5_PM_CAP_VER_ID = 3'h3;
  parameter VF5_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF5_TPHR_CAP_ENABLE = "FALSE";
  parameter VF5_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF5_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF5_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF5_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF5_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF5_TPHR_CAP_VER = 4'h1;
  
  localparam in_delay = 0;
  localparam out_delay = 0;
  localparam INCLK_DELAY = 0;
  localparam OUTCLK_DELAY = 0;

  output CFGERRCOROUT;
  output CFGERRFATALOUT;
  output CFGERRNONFATALOUT;
  output CFGEXTREADRECEIVED;
  output CFGEXTWRITERECEIVED;
  output CFGHOTRESETOUT;
  output CFGINPUTUPDATEDONE;
  output CFGINTERRUPTAOUTPUT;
  output CFGINTERRUPTBOUTPUT;
  output CFGINTERRUPTCOUTPUT;
  output CFGINTERRUPTDOUTPUT;
  output CFGINTERRUPTMSIFAIL;
  output CFGINTERRUPTMSIMASKUPDATE;
  output CFGINTERRUPTMSISENT;
  output CFGINTERRUPTMSIXFAIL;
  output CFGINTERRUPTMSIXSENT;
  output CFGINTERRUPTSENT;
  output CFGLOCALERROR;
  output CFGLTRENABLE;
  output CFGMCUPDATEDONE;
  output CFGMGMTREADWRITEDONE;
  output CFGMSGRECEIVED;
  output CFGMSGTRANSMITDONE;
  output CFGPERFUNCTIONUPDATEDONE;
  output CFGPHYLINKDOWN;
  output CFGPLSTATUSCHANGE;
  output CFGPOWERSTATECHANGEINTERRUPT;
  output CFGTPHSTTREADENABLE;
  output CFGTPHSTTWRITEENABLE;
  output DRPRDY;
  output MAXISCQTLAST;
  output MAXISCQTVALID;
  output MAXISRCTLAST;
  output MAXISRCTVALID;
  output PCIERQSEQNUMVLD;
  output PCIERQTAGVLD;
  output PIPERX0POLARITY;
  output PIPERX1POLARITY;
  output PIPERX2POLARITY;
  output PIPERX3POLARITY;
  output PIPERX4POLARITY;
  output PIPERX5POLARITY;
  output PIPERX6POLARITY;
  output PIPERX7POLARITY;
  output PIPETX0COMPLIANCE;
  output PIPETX0DATAVALID;
  output PIPETX0ELECIDLE;
  output PIPETX0STARTBLOCK;
  output PIPETX1COMPLIANCE;
  output PIPETX1DATAVALID;
  output PIPETX1ELECIDLE;
  output PIPETX1STARTBLOCK;
  output PIPETX2COMPLIANCE;
  output PIPETX2DATAVALID;
  output PIPETX2ELECIDLE;
  output PIPETX2STARTBLOCK;
  output PIPETX3COMPLIANCE;
  output PIPETX3DATAVALID;
  output PIPETX3ELECIDLE;
  output PIPETX3STARTBLOCK;
  output PIPETX4COMPLIANCE;
  output PIPETX4DATAVALID;
  output PIPETX4ELECIDLE;
  output PIPETX4STARTBLOCK;
  output PIPETX5COMPLIANCE;
  output PIPETX5DATAVALID;
  output PIPETX5ELECIDLE;
  output PIPETX5STARTBLOCK;
  output PIPETX6COMPLIANCE;
  output PIPETX6DATAVALID;
  output PIPETX6ELECIDLE;
  output PIPETX6STARTBLOCK;
  output PIPETX7COMPLIANCE;
  output PIPETX7DATAVALID;
  output PIPETX7ELECIDLE;
  output PIPETX7STARTBLOCK;
  output PIPETXDEEMPH;
  output PIPETXRCVRDET;
  output PIPETXRESET;
  output PIPETXSWING;
  output PLEQINPROGRESS;
  output [11:0] CFGFCCPLD;
  output [11:0] CFGFCNPD;
  output [11:0] CFGFCPD;
  output [11:0] CFGVFSTATUS;
  output [143:0] MIREPLAYRAMWRITEDATA;
  output [143:0] MIREQUESTRAMWRITEDATA;
  output [15:0] CFGPERFUNCSTATUSDATA;
  output [15:0] DBGDATAOUT;
  output [15:0] DRPDO;
  output [17:0] CFGVFPOWERSTATE;
  output [17:0] CFGVFTPHSTMODE;
  output [1:0] CFGDPASUBSTATECHANGE;
  output [1:0] CFGFLRINPROCESS;
  output [1:0] CFGINTERRUPTMSIENABLE;
  output [1:0] CFGINTERRUPTMSIXENABLE;
  output [1:0] CFGINTERRUPTMSIXMASK;
  output [1:0] CFGLINKPOWERSTATE;
  output [1:0] CFGOBFFENABLE;
  output [1:0] CFGPHYLINKSTATUS;
  output [1:0] CFGRCBSTATUS;
  output [1:0] CFGTPHREQUESTERENABLE;
  output [1:0] MIREPLAYRAMREADENABLE;
  output [1:0] MIREPLAYRAMWRITEENABLE;
  output [1:0] PCIERQTAGAV;
  output [1:0] PCIETFCNPDAV;
  output [1:0] PCIETFCNPHAV;
  output [1:0] PIPERX0EQCONTROL;
  output [1:0] PIPERX1EQCONTROL;
  output [1:0] PIPERX2EQCONTROL;
  output [1:0] PIPERX3EQCONTROL;
  output [1:0] PIPERX4EQCONTROL;
  output [1:0] PIPERX5EQCONTROL;
  output [1:0] PIPERX6EQCONTROL;
  output [1:0] PIPERX7EQCONTROL;
  output [1:0] PIPETX0CHARISK;
  output [1:0] PIPETX0EQCONTROL;
  output [1:0] PIPETX0POWERDOWN;
  output [1:0] PIPETX0SYNCHEADER;
  output [1:0] PIPETX1CHARISK;
  output [1:0] PIPETX1EQCONTROL;
  output [1:0] PIPETX1POWERDOWN;
  output [1:0] PIPETX1SYNCHEADER;
  output [1:0] PIPETX2CHARISK;
  output [1:0] PIPETX2EQCONTROL;
  output [1:0] PIPETX2POWERDOWN;
  output [1:0] PIPETX2SYNCHEADER;
  output [1:0] PIPETX3CHARISK;
  output [1:0] PIPETX3EQCONTROL;
  output [1:0] PIPETX3POWERDOWN;
  output [1:0] PIPETX3SYNCHEADER;
  output [1:0] PIPETX4CHARISK;
  output [1:0] PIPETX4EQCONTROL;
  output [1:0] PIPETX4POWERDOWN;
  output [1:0] PIPETX4SYNCHEADER;
  output [1:0] PIPETX5CHARISK;
  output [1:0] PIPETX5EQCONTROL;
  output [1:0] PIPETX5POWERDOWN;
  output [1:0] PIPETX5SYNCHEADER;
  output [1:0] PIPETX6CHARISK;
  output [1:0] PIPETX6EQCONTROL;
  output [1:0] PIPETX6POWERDOWN;
  output [1:0] PIPETX6SYNCHEADER;
  output [1:0] PIPETX7CHARISK;
  output [1:0] PIPETX7EQCONTROL;
  output [1:0] PIPETX7POWERDOWN;
  output [1:0] PIPETX7SYNCHEADER;
  output [1:0] PIPETXRATE;
  output [1:0] PLEQPHASE;
  output [255:0] MAXISCQTDATA;
  output [255:0] MAXISRCTDATA;
  output [2:0] CFGCURRENTSPEED;
  output [2:0] CFGMAXPAYLOAD;
  output [2:0] CFGMAXREADREQ;
  output [2:0] CFGTPHFUNCTIONNUM;
  output [2:0] PIPERX0EQPRESET;
  output [2:0] PIPERX1EQPRESET;
  output [2:0] PIPERX2EQPRESET;
  output [2:0] PIPERX3EQPRESET;
  output [2:0] PIPERX4EQPRESET;
  output [2:0] PIPERX5EQPRESET;
  output [2:0] PIPERX6EQPRESET;
  output [2:0] PIPERX7EQPRESET;
  output [2:0] PIPETXMARGIN;
  output [31:0] CFGEXTWRITEDATA;
  output [31:0] CFGINTERRUPTMSIDATA;
  output [31:0] CFGMGMTREADDATA;
  output [31:0] CFGTPHSTTWRITEDATA;
  output [31:0] PIPETX0DATA;
  output [31:0] PIPETX1DATA;
  output [31:0] PIPETX2DATA;
  output [31:0] PIPETX3DATA;
  output [31:0] PIPETX4DATA;
  output [31:0] PIPETX5DATA;
  output [31:0] PIPETX6DATA;
  output [31:0] PIPETX7DATA;
  output [3:0] CFGEXTWRITEBYTEENABLE;
  output [3:0] CFGNEGOTIATEDWIDTH;
  output [3:0] CFGTPHSTTWRITEBYTEVALID;
  output [3:0] MICOMPLETIONRAMREADENABLEL;
  output [3:0] MICOMPLETIONRAMREADENABLEU;
  output [3:0] MICOMPLETIONRAMWRITEENABLEL;
  output [3:0] MICOMPLETIONRAMWRITEENABLEU;
  output [3:0] MIREQUESTRAMREADENABLE;
  output [3:0] MIREQUESTRAMWRITEENABLE;
  output [3:0] PCIERQSEQNUM;
  output [3:0] PIPERX0EQLPTXPRESET;
  output [3:0] PIPERX1EQLPTXPRESET;
  output [3:0] PIPERX2EQLPTXPRESET;
  output [3:0] PIPERX3EQLPTXPRESET;
  output [3:0] PIPERX4EQLPTXPRESET;
  output [3:0] PIPERX5EQLPTXPRESET;
  output [3:0] PIPERX6EQLPTXPRESET;
  output [3:0] PIPERX7EQLPTXPRESET;
  output [3:0] PIPETX0EQPRESET;
  output [3:0] PIPETX1EQPRESET;
  output [3:0] PIPETX2EQPRESET;
  output [3:0] PIPETX3EQPRESET;
  output [3:0] PIPETX4EQPRESET;
  output [3:0] PIPETX5EQPRESET;
  output [3:0] PIPETX6EQPRESET;
  output [3:0] PIPETX7EQPRESET;
  output [3:0] SAXISCCTREADY;
  output [3:0] SAXISRQTREADY;
  output [4:0] CFGMSGRECEIVEDTYPE;
  output [4:0] CFGTPHSTTADDRESS;
  output [5:0] CFGFUNCTIONPOWERSTATE;
  output [5:0] CFGINTERRUPTMSIMMENABLE;
  output [5:0] CFGINTERRUPTMSIVFENABLE;
  output [5:0] CFGINTERRUPTMSIXVFENABLE;
  output [5:0] CFGINTERRUPTMSIXVFMASK;
  output [5:0] CFGLTSSMSTATE;
  output [5:0] CFGTPHSTMODE;
  output [5:0] CFGVFFLRINPROCESS;
  output [5:0] CFGVFTPHREQUESTERENABLE;
  output [5:0] PCIECQNPREQCOUNT;
  output [5:0] PCIERQTAG;
  output [5:0] PIPERX0EQLPLFFS;
  output [5:0] PIPERX1EQLPLFFS;
  output [5:0] PIPERX2EQLPLFFS;
  output [5:0] PIPERX3EQLPLFFS;
  output [5:0] PIPERX4EQLPLFFS;
  output [5:0] PIPERX5EQLPLFFS;
  output [5:0] PIPERX6EQLPLFFS;
  output [5:0] PIPERX7EQLPLFFS;
  output [5:0] PIPETX0EQDEEMPH;
  output [5:0] PIPETX1EQDEEMPH;
  output [5:0] PIPETX2EQDEEMPH;
  output [5:0] PIPETX3EQDEEMPH;
  output [5:0] PIPETX4EQDEEMPH;
  output [5:0] PIPETX5EQDEEMPH;
  output [5:0] PIPETX6EQDEEMPH;
  output [5:0] PIPETX7EQDEEMPH;
  output [71:0] MICOMPLETIONRAMWRITEDATAL;
  output [71:0] MICOMPLETIONRAMWRITEDATAU;
  output [74:0] MAXISRCTUSER;
  output [7:0] CFGEXTFUNCTIONNUMBER;
  output [7:0] CFGFCCPLH;
  output [7:0] CFGFCNPH;
  output [7:0] CFGFCPH;
  output [7:0] CFGFUNCTIONSTATUS;
  output [7:0] CFGMSGRECEIVEDDATA;
  output [7:0] MAXISCQTKEEP;
  output [7:0] MAXISRCTKEEP;
  output [7:0] PLGEN3PCSRXSLIDE;
  output [84:0] MAXISCQTUSER;
  output [8:0] MIREPLAYRAMADDRESS;
  output [8:0] MIREQUESTRAMREADADDRESSA;
  output [8:0] MIREQUESTRAMREADADDRESSB;
  output [8:0] MIREQUESTRAMWRITEADDRESSA;
  output [8:0] MIREQUESTRAMWRITEADDRESSB;
  output [9:0] CFGEXTREGISTERNUMBER;
  output [9:0] MICOMPLETIONRAMREADADDRESSAL;
  output [9:0] MICOMPLETIONRAMREADADDRESSAU;
  output [9:0] MICOMPLETIONRAMREADADDRESSBL;
  output [9:0] MICOMPLETIONRAMREADADDRESSBU;
  output [9:0] MICOMPLETIONRAMWRITEADDRESSAL;
  output [9:0] MICOMPLETIONRAMWRITEADDRESSAU;
  output [9:0] MICOMPLETIONRAMWRITEADDRESSBL;
  output [9:0] MICOMPLETIONRAMWRITEADDRESSBU;

  input CFGCONFIGSPACEENABLE;
  input CFGERRCORIN;
  input CFGERRUNCORIN;
  input CFGEXTREADDATAVALID;
  input CFGHOTRESETIN;
  input CFGINPUTUPDATEREQUEST;
  input CFGINTERRUPTMSITPHPRESENT;
  input CFGINTERRUPTMSIXINT;
  input CFGLINKTRAININGENABLE;
  input CFGMCUPDATEREQUEST;
  input CFGMGMTREAD;
  input CFGMGMTTYPE1CFGREGACCESS;
  input CFGMGMTWRITE;
  input CFGMSGTRANSMIT;
  input CFGPERFUNCTIONOUTPUTREQUEST;
  input CFGPOWERSTATECHANGEACK;
  input CFGREQPMTRANSITIONL23READY;
  input CFGTPHSTTREADDATAVALID;
  input CORECLK;
  input CORECLKMICOMPLETIONRAML;
  input CORECLKMICOMPLETIONRAMU;
  input CORECLKMIREPLAYRAM;
  input CORECLKMIREQUESTRAM;
  input DRPCLK;
  input DRPEN;
  input DRPWE;
  input MGMTRESETN;
  input MGMTSTICKYRESETN;
  input PCIECQNPREQ;
  input PIPECLK;
  input PIPERESETN;
  input PIPERX0DATAVALID;
  input PIPERX0ELECIDLE;
  input PIPERX0EQDONE;
  input PIPERX0EQLPADAPTDONE;
  input PIPERX0EQLPLFFSSEL;
  input PIPERX0PHYSTATUS;
  input PIPERX0STARTBLOCK;
  input PIPERX0VALID;
  input PIPERX1DATAVALID;
  input PIPERX1ELECIDLE;
  input PIPERX1EQDONE;
  input PIPERX1EQLPADAPTDONE;
  input PIPERX1EQLPLFFSSEL;
  input PIPERX1PHYSTATUS;
  input PIPERX1STARTBLOCK;
  input PIPERX1VALID;
  input PIPERX2DATAVALID;
  input PIPERX2ELECIDLE;
  input PIPERX2EQDONE;
  input PIPERX2EQLPADAPTDONE;
  input PIPERX2EQLPLFFSSEL;
  input PIPERX2PHYSTATUS;
  input PIPERX2STARTBLOCK;
  input PIPERX2VALID;
  input PIPERX3DATAVALID;
  input PIPERX3ELECIDLE;
  input PIPERX3EQDONE;
  input PIPERX3EQLPADAPTDONE;
  input PIPERX3EQLPLFFSSEL;
  input PIPERX3PHYSTATUS;
  input PIPERX3STARTBLOCK;
  input PIPERX3VALID;
  input PIPERX4DATAVALID;
  input PIPERX4ELECIDLE;
  input PIPERX4EQDONE;
  input PIPERX4EQLPADAPTDONE;
  input PIPERX4EQLPLFFSSEL;
  input PIPERX4PHYSTATUS;
  input PIPERX4STARTBLOCK;
  input PIPERX4VALID;
  input PIPERX5DATAVALID;
  input PIPERX5ELECIDLE;
  input PIPERX5EQDONE;
  input PIPERX5EQLPADAPTDONE;
  input PIPERX5EQLPLFFSSEL;
  input PIPERX5PHYSTATUS;
  input PIPERX5STARTBLOCK;
  input PIPERX5VALID;
  input PIPERX6DATAVALID;
  input PIPERX6ELECIDLE;
  input PIPERX6EQDONE;
  input PIPERX6EQLPADAPTDONE;
  input PIPERX6EQLPLFFSSEL;
  input PIPERX6PHYSTATUS;
  input PIPERX6STARTBLOCK;
  input PIPERX6VALID;
  input PIPERX7DATAVALID;
  input PIPERX7ELECIDLE;
  input PIPERX7EQDONE;
  input PIPERX7EQLPADAPTDONE;
  input PIPERX7EQLPLFFSSEL;
  input PIPERX7PHYSTATUS;
  input PIPERX7STARTBLOCK;
  input PIPERX7VALID;
  input PIPETX0EQDONE;
  input PIPETX1EQDONE;
  input PIPETX2EQDONE;
  input PIPETX3EQDONE;
  input PIPETX4EQDONE;
  input PIPETX5EQDONE;
  input PIPETX6EQDONE;
  input PIPETX7EQDONE;
  input PLDISABLESCRAMBLER;
  input PLEQRESETEIEOSCOUNT;
  input PLGEN3PCSDISABLE;
  input RECCLK;
  input RESETN;
  input SAXISCCTLAST;
  input SAXISCCTVALID;
  input SAXISRQTLAST;
  input SAXISRQTVALID;
  input USERCLK;
  input [10:0] DRPADDR;
  input [143:0] MICOMPLETIONRAMREADDATA;
  input [143:0] MIREPLAYRAMREADDATA;
  input [143:0] MIREQUESTRAMREADDATA;
  input [15:0] CFGDEVID;
  input [15:0] CFGSUBSYSID;
  input [15:0] CFGSUBSYSVENDID;
  input [15:0] CFGVENDID;
  input [15:0] DRPDI;
  input [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPETX0EQCOEFF;
  input [17:0] PIPETX1EQCOEFF;
  input [17:0] PIPETX2EQCOEFF;
  input [17:0] PIPETX3EQCOEFF;
  input [17:0] PIPETX4EQCOEFF;
  input [17:0] PIPETX5EQCOEFF;
  input [17:0] PIPETX6EQCOEFF;
  input [17:0] PIPETX7EQCOEFF;
  input [18:0] CFGMGMTADDR;
  input [1:0] CFGFLRDONE;
  input [1:0] CFGINTERRUPTMSITPHTYPE;
  input [1:0] CFGINTERRUPTPENDING;
  input [1:0] PIPERX0CHARISK;
  input [1:0] PIPERX0SYNCHEADER;
  input [1:0] PIPERX1CHARISK;
  input [1:0] PIPERX1SYNCHEADER;
  input [1:0] PIPERX2CHARISK;
  input [1:0] PIPERX2SYNCHEADER;
  input [1:0] PIPERX3CHARISK;
  input [1:0] PIPERX3SYNCHEADER;
  input [1:0] PIPERX4CHARISK;
  input [1:0] PIPERX4SYNCHEADER;
  input [1:0] PIPERX5CHARISK;
  input [1:0] PIPERX5SYNCHEADER;
  input [1:0] PIPERX6CHARISK;
  input [1:0] PIPERX6SYNCHEADER;
  input [1:0] PIPERX7CHARISK;
  input [1:0] PIPERX7SYNCHEADER;
  input [21:0] MAXISCQTREADY;
  input [21:0] MAXISRCTREADY;
  input [255:0] SAXISCCTDATA;
  input [255:0] SAXISRQTDATA;
  input [2:0] CFGDSFUNCTIONNUMBER;
  input [2:0] CFGFCSEL;
  input [2:0] CFGINTERRUPTMSIATTR;
  input [2:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
  input [2:0] CFGMSGTRANSMITTYPE;
  input [2:0] CFGPERFUNCSTATUSCONTROL;
  input [2:0] CFGPERFUNCTIONNUMBER;
  input [2:0] PIPERX0STATUS;
  input [2:0] PIPERX1STATUS;
  input [2:0] PIPERX2STATUS;
  input [2:0] PIPERX3STATUS;
  input [2:0] PIPERX4STATUS;
  input [2:0] PIPERX5STATUS;
  input [2:0] PIPERX6STATUS;
  input [2:0] PIPERX7STATUS;
  input [31:0] CFGEXTREADDATA;
  input [31:0] CFGINTERRUPTMSIINT;
  input [31:0] CFGINTERRUPTMSIXDATA;
  input [31:0] CFGMGMTWRITEDATA;
  input [31:0] CFGMSGTRANSMITDATA;
  input [31:0] CFGTPHSTTREADDATA;
  input [31:0] PIPERX0DATA;
  input [31:0] PIPERX1DATA;
  input [31:0] PIPERX2DATA;
  input [31:0] PIPERX3DATA;
  input [31:0] PIPERX4DATA;
  input [31:0] PIPERX5DATA;
  input [31:0] PIPERX6DATA;
  input [31:0] PIPERX7DATA;
  input [32:0] SAXISCCTUSER;
  input [3:0] CFGINTERRUPTINT;
  input [3:0] CFGINTERRUPTMSISELECT;
  input [3:0] CFGMGMTBYTEENABLE;
  input [4:0] CFGDSDEVICENUMBER;
  input [59:0] SAXISRQTUSER;
  input [5:0] CFGVFFLRDONE;
  input [5:0] PIPEEQFS;
  input [5:0] PIPEEQLF;
  input [63:0] CFGDSN;
  input [63:0] CFGINTERRUPTMSIPENDINGSTATUS;
  input [63:0] CFGINTERRUPTMSIXADDRESS;
  input [7:0] CFGDSBUSNUMBER;
  input [7:0] CFGDSPORTNUMBER;
  input [7:0] CFGREVID;
  input [7:0] PLGEN3PCSRXSYNCDONE;
  input [7:0] SAXISCCTKEEP;
  input [7:0] SAXISRQTKEEP;
  input [8:0] CFGINTERRUPTMSITPHSTTAG;

  reg SIM_VERSION_BINARY;
  reg [0:0] ARI_CAP_ENABLE_BINARY;
  reg [0:0] AXISTEN_IF_CC_ALIGNMENT_MODE_BINARY;
  reg [0:0] AXISTEN_IF_CC_PARITY_CHK_BINARY;
  reg [0:0] AXISTEN_IF_CQ_ALIGNMENT_MODE_BINARY;
  reg [0:0] AXISTEN_IF_ENABLE_CLIENT_TAG_BINARY;
  reg [0:0] AXISTEN_IF_ENABLE_RX_MSG_INTFC_BINARY;
  reg [0:0] AXISTEN_IF_RC_ALIGNMENT_MODE_BINARY;
  reg [0:0] AXISTEN_IF_RC_STRADDLE_BINARY;
  reg [0:0] AXISTEN_IF_RQ_ALIGNMENT_MODE_BINARY;
  reg [0:0] AXISTEN_IF_RQ_PARITY_CHK_BINARY;
  reg [0:0] CRM_CORE_CLK_FREQ_500_BINARY;
  reg [0:0] GEN3_PCS_RX_ELECIDLE_INTERNAL_BINARY;
  reg [0:0] LL_ACK_TIMEOUT_EN_BINARY;
  reg [0:0] LL_CPL_FC_UPDATE_TIMER_OVERRIDE_BINARY;
  reg [0:0] LL_FC_UPDATE_TIMER_OVERRIDE_BINARY;
  reg [0:0] LL_NP_FC_UPDATE_TIMER_OVERRIDE_BINARY;
  reg [0:0] LL_P_FC_UPDATE_TIMER_OVERRIDE_BINARY;
  reg [0:0] LL_REPLAY_TIMEOUT_EN_BINARY;
  reg [0:0] LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_BINARY;
  reg [0:0] LTR_TX_MESSAGE_ON_LTR_ENABLE_BINARY;
  reg [0:0] PF0_AER_CAP_ECRC_CHECK_CAPABLE_BINARY;
  reg [0:0] PF0_AER_CAP_ECRC_GEN_CAPABLE_BINARY;
  reg [0:0] PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_BINARY;
  reg [0:0] PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_BINARY;
  reg [0:0] PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_BINARY;
  reg [0:0] PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_BINARY;
  reg [0:0] PF0_DEV_CAP2_LTR_SUPPORT_BINARY;
  reg [0:0] PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_BINARY;
  reg [0:0] PF0_DEV_CAP_EXT_TAG_SUPPORTED_BINARY;
  reg [0:0] PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_BINARY;
  reg [0:0] PF0_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY;
  reg [0:0] PF0_EXPANSION_ROM_ENABLE_BINARY;
  reg [0:0] PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_BINARY;
  reg [0:0] PF0_PB_CAP_SYSTEM_ALLOCATED_BINARY;
  reg [0:0] PF0_PM_CAP_PMESUPPORT_D0_BINARY;
  reg [0:0] PF0_PM_CAP_PMESUPPORT_D1_BINARY;
  reg [0:0] PF0_PM_CAP_PMESUPPORT_D3HOT_BINARY;
  reg [0:0] PF0_PM_CAP_SUPP_D1_STATE_BINARY;
  reg [0:0] PF0_PM_CSR_NOSOFTRESET_BINARY;
  reg [0:0] PF0_RBAR_CAP_ENABLE_BINARY;
  reg [0:0] PF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] PF0_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] PF0_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] PF1_AER_CAP_ECRC_CHECK_CAPABLE_BINARY;
  reg [0:0] PF1_AER_CAP_ECRC_GEN_CAPABLE_BINARY;
  reg [0:0] PF1_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY;
  reg [0:0] PF1_EXPANSION_ROM_ENABLE_BINARY;
  reg [0:0] PF1_PB_CAP_SYSTEM_ALLOCATED_BINARY;
  reg [0:0] PF1_RBAR_CAP_ENABLE_BINARY;
  reg [0:0] PF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] PF1_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] PF1_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] PL_DISABLE_EI_INFER_IN_L0_BINARY;
  reg [0:0] PL_DISABLE_GEN3_DC_BALANCE_BINARY;
  reg [0:0] PL_DISABLE_SCRAMBLING_BINARY;
  reg [0:0] PL_DISABLE_UPCONFIG_CAPABLE_BINARY;
  reg [0:0] PL_EQ_ADAPT_DISABLE_COEFF_CHECK_BINARY;
  reg [0:0] PL_EQ_ADAPT_DISABLE_PRESET_CHECK_BINARY;
  reg [0:0] PL_EQ_BYPASS_PHASE23_BINARY;
  reg [0:0] PL_EQ_SHORT_ADAPT_PHASE_BINARY;
  reg [0:0] PL_SIM_FAST_LINK_TRAINING_BINARY;
  reg [0:0] PL_UPSTREAM_FACING_BINARY;
  reg [0:0] PM_ENABLE_SLOT_POWER_CAPTURE_BINARY;
  reg [0:0] SPARE_BIT0_BINARY;
  reg [0:0] SPARE_BIT1_BINARY;
  reg [0:0] SPARE_BIT2_BINARY;
  reg [0:0] SPARE_BIT3_BINARY;
  reg [0:0] SPARE_BIT4_BINARY;
  reg [0:0] SPARE_BIT5_BINARY;
  reg [0:0] SPARE_BIT6_BINARY;
  reg [0:0] SPARE_BIT7_BINARY;
  reg [0:0] SPARE_BIT8_BINARY;
  reg [0:0] SRIOV_CAP_ENABLE_BINARY;
  reg [0:0] TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_BINARY;
  reg [0:0] TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_BINARY;
  reg [0:0] TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_BINARY;
  reg [0:0] TL_LEGACY_MODE_ENABLE_BINARY;
  reg [0:0] TL_PF_ENABLE_REG_BINARY;
  reg [0:0] TL_TAG_MGMT_ENABLE_BINARY;
  reg [0:0] VF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF0_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF0_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] VF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF1_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF1_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] VF2_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF2_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF2_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] VF3_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF3_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF3_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] VF4_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF4_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF4_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] VF5_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF5_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF5_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [1:0] LL_ACK_TIMEOUT_FUNC_BINARY;
  reg [1:0] LL_REPLAY_TIMEOUT_FUNC_BINARY;
  reg [1:0] PF0_LINK_CAP_ASPM_SUPPORT_BINARY;
  reg [2:0] PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_BINARY;
  reg [2:0] PF0_DEV_CAP_ENDPOINT_L1_LATENCY_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_BINARY;
  reg [2:0] PF0_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] PF0_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] PF0_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] PF1_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] PF1_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] PF1_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF0_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF0_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF0_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF1_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF1_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF1_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF2_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF2_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF2_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF3_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF3_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF3_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF4_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF4_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF4_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF5_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF5_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF5_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [7:0] PL_N_FTS_COMCLK_GEN1_BINARY;
  reg [7:0] PL_N_FTS_COMCLK_GEN2_BINARY;
  reg [7:0] PL_N_FTS_COMCLK_GEN3_BINARY;
  reg [7:0] PL_N_FTS_GEN1_BINARY;
  reg [7:0] PL_N_FTS_GEN2_BINARY;
  reg [7:0] PL_N_FTS_GEN3_BINARY;

  reg notifier;

  initial begin
    case (ARI_CAP_ENABLE)
      "FALSE" : ARI_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : ARI_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute ARI_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", ARI_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (AXISTEN_IF_CC_ALIGNMENT_MODE)
      "FALSE" : AXISTEN_IF_CC_ALIGNMENT_MODE_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_CC_ALIGNMENT_MODE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_CC_ALIGNMENT_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_CC_ALIGNMENT_MODE);
        #1 $finish;
      end
    endcase

    case (AXISTEN_IF_CC_PARITY_CHK)
      "TRUE" : AXISTEN_IF_CC_PARITY_CHK_BINARY = 1'b1;
      "FALSE" : AXISTEN_IF_CC_PARITY_CHK_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_CC_PARITY_CHK on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", AXISTEN_IF_CC_PARITY_CHK);
        #1 $finish;
      end
    endcase

    case (AXISTEN_IF_CQ_ALIGNMENT_MODE)
      "FALSE" : AXISTEN_IF_CQ_ALIGNMENT_MODE_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_CQ_ALIGNMENT_MODE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_CQ_ALIGNMENT_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_CQ_ALIGNMENT_MODE);
        #1 $finish;
      end
    endcase

    case (AXISTEN_IF_ENABLE_CLIENT_TAG)
      "FALSE" : AXISTEN_IF_ENABLE_CLIENT_TAG_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_ENABLE_CLIENT_TAG_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_ENABLE_CLIENT_TAG on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_ENABLE_CLIENT_TAG);
        #1 $finish;
      end
    endcase

    case (AXISTEN_IF_ENABLE_RX_MSG_INTFC)
      "FALSE" : AXISTEN_IF_ENABLE_RX_MSG_INTFC_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_ENABLE_RX_MSG_INTFC_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_ENABLE_RX_MSG_INTFC on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_ENABLE_RX_MSG_INTFC);
        #1 $finish;
      end
    endcase

    case (AXISTEN_IF_RC_ALIGNMENT_MODE)
      "FALSE" : AXISTEN_IF_RC_ALIGNMENT_MODE_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_RC_ALIGNMENT_MODE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_RC_ALIGNMENT_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_RC_ALIGNMENT_MODE);
        #1 $finish;
      end
    endcase

    case (AXISTEN_IF_RC_STRADDLE)
      "FALSE" : AXISTEN_IF_RC_STRADDLE_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_RC_STRADDLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_RC_STRADDLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_RC_STRADDLE);
        #1 $finish;
      end
    endcase

    case (AXISTEN_IF_RQ_ALIGNMENT_MODE)
      "FALSE" : AXISTEN_IF_RQ_ALIGNMENT_MODE_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_RQ_ALIGNMENT_MODE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_RQ_ALIGNMENT_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_RQ_ALIGNMENT_MODE);
        #1 $finish;
      end
    endcase

    case (AXISTEN_IF_RQ_PARITY_CHK)
      "TRUE" : AXISTEN_IF_RQ_PARITY_CHK_BINARY = 1'b1;
      "FALSE" : AXISTEN_IF_RQ_PARITY_CHK_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_RQ_PARITY_CHK on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", AXISTEN_IF_RQ_PARITY_CHK);
        #1 $finish;
      end
    endcase

    case (CRM_CORE_CLK_FREQ_500)
      "TRUE" : CRM_CORE_CLK_FREQ_500_BINARY = 1'b1;
      "FALSE" : CRM_CORE_CLK_FREQ_500_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute CRM_CORE_CLK_FREQ_500 on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", CRM_CORE_CLK_FREQ_500);
        #1 $finish;
      end
    endcase

    case (GEN3_PCS_RX_ELECIDLE_INTERNAL)
      "TRUE" : GEN3_PCS_RX_ELECIDLE_INTERNAL_BINARY = 1'b1;
      "FALSE" : GEN3_PCS_RX_ELECIDLE_INTERNAL_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute GEN3_PCS_RX_ELECIDLE_INTERNAL on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", GEN3_PCS_RX_ELECIDLE_INTERNAL);
        #1 $finish;
      end
    endcase

    case (LL_ACK_TIMEOUT_EN)
      "FALSE" : LL_ACK_TIMEOUT_EN_BINARY = 1'b0;
      "TRUE" : LL_ACK_TIMEOUT_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_ACK_TIMEOUT_EN on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_ACK_TIMEOUT_EN);
        #1 $finish;
      end
    endcase

    case (LL_CPL_FC_UPDATE_TIMER_OVERRIDE)
      "FALSE" : LL_CPL_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b0;
      "TRUE" : LL_CPL_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_CPL_FC_UPDATE_TIMER_OVERRIDE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_CPL_FC_UPDATE_TIMER_OVERRIDE);
        #1 $finish;
      end
    endcase

    case (LL_FC_UPDATE_TIMER_OVERRIDE)
      "FALSE" : LL_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b0;
      "TRUE" : LL_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_FC_UPDATE_TIMER_OVERRIDE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_FC_UPDATE_TIMER_OVERRIDE);
        #1 $finish;
      end
    endcase

    case (LL_NP_FC_UPDATE_TIMER_OVERRIDE)
      "FALSE" : LL_NP_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b0;
      "TRUE" : LL_NP_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_NP_FC_UPDATE_TIMER_OVERRIDE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_NP_FC_UPDATE_TIMER_OVERRIDE);
        #1 $finish;
      end
    endcase

    case (LL_P_FC_UPDATE_TIMER_OVERRIDE)
      "FALSE" : LL_P_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b0;
      "TRUE" : LL_P_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_P_FC_UPDATE_TIMER_OVERRIDE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_P_FC_UPDATE_TIMER_OVERRIDE);
        #1 $finish;
      end
    endcase

    case (LL_REPLAY_TIMEOUT_EN)
      "FALSE" : LL_REPLAY_TIMEOUT_EN_BINARY = 1'b0;
      "TRUE" : LL_REPLAY_TIMEOUT_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_REPLAY_TIMEOUT_EN on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_REPLAY_TIMEOUT_EN);
        #1 $finish;
      end
    endcase

    case (LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE)
      "FALSE" : LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_BINARY = 1'b0;
      "TRUE" : LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE);
        #1 $finish;
      end
    endcase

    case (LTR_TX_MESSAGE_ON_LTR_ENABLE)
      "FALSE" : LTR_TX_MESSAGE_ON_LTR_ENABLE_BINARY = 1'b0;
      "TRUE" : LTR_TX_MESSAGE_ON_LTR_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LTR_TX_MESSAGE_ON_LTR_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LTR_TX_MESSAGE_ON_LTR_ENABLE);
        #1 $finish;
      end
    endcase

    case (PF0_AER_CAP_ECRC_CHECK_CAPABLE)
      "FALSE" : PF0_AER_CAP_ECRC_CHECK_CAPABLE_BINARY = 1'b0;
      "TRUE" : PF0_AER_CAP_ECRC_CHECK_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_AER_CAP_ECRC_CHECK_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_AER_CAP_ECRC_CHECK_CAPABLE);
        #1 $finish;
      end
    endcase

    case (PF0_AER_CAP_ECRC_GEN_CAPABLE)
      "FALSE" : PF0_AER_CAP_ECRC_GEN_CAPABLE_BINARY = 1'b0;
      "TRUE" : PF0_AER_CAP_ECRC_GEN_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_AER_CAP_ECRC_GEN_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_AER_CAP_ECRC_GEN_CAPABLE);
        #1 $finish;
      end
    endcase

    case (PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT)
      "TRUE" : PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT);
        #1 $finish;
      end
    endcase

    case (PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT)
      "TRUE" : PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT);
        #1 $finish;
      end
    endcase

    case (PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT)
      "TRUE" : PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT);
        #1 $finish;
      end
    endcase

    case (PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE)
      "TRUE" : PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE);
        #1 $finish;
      end
    endcase

    case (PF0_DEV_CAP2_LTR_SUPPORT)
      "TRUE" : PF0_DEV_CAP2_LTR_SUPPORT_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP2_LTR_SUPPORT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_LTR_SUPPORT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP2_LTR_SUPPORT);
        #1 $finish;
      end
    endcase

    case (PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT)
      "FALSE" : PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_BINARY = 1'b0;
      "TRUE" : PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT);
        #1 $finish;
      end
    endcase

    case (PF0_DEV_CAP_EXT_TAG_SUPPORTED)
      "TRUE" : PF0_DEV_CAP_EXT_TAG_SUPPORTED_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP_EXT_TAG_SUPPORTED_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP_EXT_TAG_SUPPORTED on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP_EXT_TAG_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE)
      "TRUE" : PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE);
        #1 $finish;
      end
    endcase

    case (PF0_DPA_CAP_SUB_STATE_CONTROL_EN)
      "TRUE" : PF0_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY = 1'b1;
      "FALSE" : PF0_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DPA_CAP_SUB_STATE_CONTROL_EN on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DPA_CAP_SUB_STATE_CONTROL_EN);
        #1 $finish;
      end
    endcase

    case (PF0_EXPANSION_ROM_ENABLE)
      "FALSE" : PF0_EXPANSION_ROM_ENABLE_BINARY = 1'b0;
      "TRUE" : PF0_EXPANSION_ROM_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_EXPANSION_ROM_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_EXPANSION_ROM_ENABLE);
        #1 $finish;
      end
    endcase

    case (PF0_LINK_STATUS_SLOT_CLOCK_CONFIG)
      "TRUE" : PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_BINARY = 1'b1;
      "FALSE" : PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_LINK_STATUS_SLOT_CLOCK_CONFIG on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_LINK_STATUS_SLOT_CLOCK_CONFIG);
        #1 $finish;
      end
    endcase

    case (PF0_PB_CAP_SYSTEM_ALLOCATED)
      "FALSE" : PF0_PB_CAP_SYSTEM_ALLOCATED_BINARY = 1'b0;
      "TRUE" : PF0_PB_CAP_SYSTEM_ALLOCATED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PB_CAP_SYSTEM_ALLOCATED on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_PB_CAP_SYSTEM_ALLOCATED);
        #1 $finish;
      end
    endcase

    case (PF0_PM_CAP_PMESUPPORT_D0)
      "TRUE" : PF0_PM_CAP_PMESUPPORT_D0_BINARY = 1'b1;
      "FALSE" : PF0_PM_CAP_PMESUPPORT_D0_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PM_CAP_PMESUPPORT_D0 on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_PM_CAP_PMESUPPORT_D0);
        #1 $finish;
      end
    endcase

    case (PF0_PM_CAP_PMESUPPORT_D1)
      "TRUE" : PF0_PM_CAP_PMESUPPORT_D1_BINARY = 1'b1;
      "FALSE" : PF0_PM_CAP_PMESUPPORT_D1_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PM_CAP_PMESUPPORT_D1 on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_PM_CAP_PMESUPPORT_D1);
        #1 $finish;
      end
    endcase

    case (PF0_PM_CAP_PMESUPPORT_D3HOT)
      "TRUE" : PF0_PM_CAP_PMESUPPORT_D3HOT_BINARY = 1'b1;
      "FALSE" : PF0_PM_CAP_PMESUPPORT_D3HOT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PM_CAP_PMESUPPORT_D3HOT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_PM_CAP_PMESUPPORT_D3HOT);
        #1 $finish;
      end
    endcase

    case (PF0_PM_CAP_SUPP_D1_STATE)
      "TRUE" : PF0_PM_CAP_SUPP_D1_STATE_BINARY = 1'b1;
      "FALSE" : PF0_PM_CAP_SUPP_D1_STATE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PM_CAP_SUPP_D1_STATE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_PM_CAP_SUPP_D1_STATE);
        #1 $finish;
      end
    endcase

    case (PF0_PM_CSR_NOSOFTRESET)
      "TRUE" : PF0_PM_CSR_NOSOFTRESET_BINARY = 1'b1;
      "FALSE" : PF0_PM_CSR_NOSOFTRESET_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PM_CSR_NOSOFTRESET on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_PM_CSR_NOSOFTRESET);
        #1 $finish;
      end
    endcase

    case (PF0_RBAR_CAP_ENABLE)
      "FALSE" : PF0_RBAR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : PF0_RBAR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_RBAR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_RBAR_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (PF0_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : PF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : PF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_TPHR_CAP_DEV_SPECIFIC_MODE);
        #1 $finish;
      end
    endcase

    case (PF0_TPHR_CAP_ENABLE)
      "FALSE" : PF0_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : PF0_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_TPHR_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (PF0_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : PF0_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : PF0_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_TPHR_CAP_INT_VEC_MODE);
        #1 $finish;
      end
    endcase

    case (PF1_AER_CAP_ECRC_CHECK_CAPABLE)
      "FALSE" : PF1_AER_CAP_ECRC_CHECK_CAPABLE_BINARY = 1'b0;
      "TRUE" : PF1_AER_CAP_ECRC_CHECK_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_AER_CAP_ECRC_CHECK_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_AER_CAP_ECRC_CHECK_CAPABLE);
        #1 $finish;
      end
    endcase

    case (PF1_AER_CAP_ECRC_GEN_CAPABLE)
      "FALSE" : PF1_AER_CAP_ECRC_GEN_CAPABLE_BINARY = 1'b0;
      "TRUE" : PF1_AER_CAP_ECRC_GEN_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_AER_CAP_ECRC_GEN_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_AER_CAP_ECRC_GEN_CAPABLE);
        #1 $finish;
      end
    endcase

    case (PF1_DPA_CAP_SUB_STATE_CONTROL_EN)
      "TRUE" : PF1_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY = 1'b1;
      "FALSE" : PF1_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_DPA_CAP_SUB_STATE_CONTROL_EN on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF1_DPA_CAP_SUB_STATE_CONTROL_EN);
        #1 $finish;
      end
    endcase

    case (PF1_EXPANSION_ROM_ENABLE)
      "FALSE" : PF1_EXPANSION_ROM_ENABLE_BINARY = 1'b0;
      "TRUE" : PF1_EXPANSION_ROM_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_EXPANSION_ROM_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_EXPANSION_ROM_ENABLE);
        #1 $finish;
      end
    endcase

    case (PF1_PB_CAP_SYSTEM_ALLOCATED)
      "FALSE" : PF1_PB_CAP_SYSTEM_ALLOCATED_BINARY = 1'b0;
      "TRUE" : PF1_PB_CAP_SYSTEM_ALLOCATED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_PB_CAP_SYSTEM_ALLOCATED on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_PB_CAP_SYSTEM_ALLOCATED);
        #1 $finish;
      end
    endcase

    case (PF1_RBAR_CAP_ENABLE)
      "FALSE" : PF1_RBAR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : PF1_RBAR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_RBAR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_RBAR_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (PF1_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : PF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : PF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF1_TPHR_CAP_DEV_SPECIFIC_MODE);
        #1 $finish;
      end
    endcase

    case (PF1_TPHR_CAP_ENABLE)
      "FALSE" : PF1_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : PF1_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_TPHR_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (PF1_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : PF1_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : PF1_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF1_TPHR_CAP_INT_VEC_MODE);
        #1 $finish;
      end
    endcase

    case (PL_DISABLE_EI_INFER_IN_L0)
      "FALSE" : PL_DISABLE_EI_INFER_IN_L0_BINARY = 1'b0;
      "TRUE" : PL_DISABLE_EI_INFER_IN_L0_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_DISABLE_EI_INFER_IN_L0 on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_DISABLE_EI_INFER_IN_L0);
        #1 $finish;
      end
    endcase

    case (PL_DISABLE_GEN3_DC_BALANCE)
      "FALSE" : PL_DISABLE_GEN3_DC_BALANCE_BINARY = 1'b0;
      "TRUE" : PL_DISABLE_GEN3_DC_BALANCE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_DISABLE_GEN3_DC_BALANCE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_DISABLE_GEN3_DC_BALANCE);
        #1 $finish;
      end
    endcase

    case (PL_DISABLE_SCRAMBLING)
      "FALSE" : PL_DISABLE_SCRAMBLING_BINARY = 1'b0;
      "TRUE" : PL_DISABLE_SCRAMBLING_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_DISABLE_SCRAMBLING on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_DISABLE_SCRAMBLING);
        #1 $finish;
      end
    endcase

    case (PL_DISABLE_UPCONFIG_CAPABLE)
      "FALSE" : PL_DISABLE_UPCONFIG_CAPABLE_BINARY = 1'b0;
      "TRUE" : PL_DISABLE_UPCONFIG_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_DISABLE_UPCONFIG_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_DISABLE_UPCONFIG_CAPABLE);
        #1 $finish;
      end
    endcase

    case (PL_EQ_ADAPT_DISABLE_COEFF_CHECK)
      "FALSE" : PL_EQ_ADAPT_DISABLE_COEFF_CHECK_BINARY = 1'b0;
      "TRUE" : PL_EQ_ADAPT_DISABLE_COEFF_CHECK_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_EQ_ADAPT_DISABLE_COEFF_CHECK on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_EQ_ADAPT_DISABLE_COEFF_CHECK);
        #1 $finish;
      end
    endcase

    case (PL_EQ_ADAPT_DISABLE_PRESET_CHECK)
      "FALSE" : PL_EQ_ADAPT_DISABLE_PRESET_CHECK_BINARY = 1'b0;
      "TRUE" : PL_EQ_ADAPT_DISABLE_PRESET_CHECK_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_EQ_ADAPT_DISABLE_PRESET_CHECK on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_EQ_ADAPT_DISABLE_PRESET_CHECK);
        #1 $finish;
      end
    endcase

    case (PL_EQ_BYPASS_PHASE23)
      "FALSE" : PL_EQ_BYPASS_PHASE23_BINARY = 1'b0;
      "TRUE" : PL_EQ_BYPASS_PHASE23_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_EQ_BYPASS_PHASE23 on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_EQ_BYPASS_PHASE23);
        #1 $finish;
      end
    endcase

    case (PL_EQ_SHORT_ADAPT_PHASE)
      "FALSE" : PL_EQ_SHORT_ADAPT_PHASE_BINARY = 1'b0;
      "TRUE" : PL_EQ_SHORT_ADAPT_PHASE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_EQ_SHORT_ADAPT_PHASE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_EQ_SHORT_ADAPT_PHASE);
        #1 $finish;
      end
    endcase

    case (PL_SIM_FAST_LINK_TRAINING)
      "FALSE" : PL_SIM_FAST_LINK_TRAINING_BINARY = 1'b0;
      "TRUE" : PL_SIM_FAST_LINK_TRAINING_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_SIM_FAST_LINK_TRAINING on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_SIM_FAST_LINK_TRAINING);
        #1 $finish;
      end
    endcase

    case (PL_UPSTREAM_FACING)
      "TRUE" : PL_UPSTREAM_FACING_BINARY = 1'b1;
      "FALSE" : PL_UPSTREAM_FACING_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_UPSTREAM_FACING on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PL_UPSTREAM_FACING);
        #1 $finish;
      end
    endcase

    case (PM_ENABLE_SLOT_POWER_CAPTURE)
      "TRUE" : PM_ENABLE_SLOT_POWER_CAPTURE_BINARY = 1'b1;
      "FALSE" : PM_ENABLE_SLOT_POWER_CAPTURE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_ENABLE_SLOT_POWER_CAPTURE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PM_ENABLE_SLOT_POWER_CAPTURE);
        #1 $finish;
      end
    endcase

    case (SIM_VERSION)
      "1.0" : SIM_VERSION_BINARY = 0;
      "1.1" : SIM_VERSION_BINARY = 0;
      "1.2" : SIM_VERSION_BINARY = 0;
      "1.3" : SIM_VERSION_BINARY = 0;
      "2.0" : SIM_VERSION_BINARY = 0;
      "3.0" : SIM_VERSION_BINARY = 0;
      "4.0" : SIM_VERSION_BINARY = 0;
      default : begin
        $display("Attribute Syntax Error : The Attribute SIM_VERSION on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are 1.0, 1.1, 1.2, 1.3, 2.0, 3.0, or 4.0.", SIM_VERSION);
        #1 $finish;
      end
    endcase

    case (SRIOV_CAP_ENABLE)
      "FALSE" : SRIOV_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : SRIOV_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SRIOV_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SRIOV_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (TL_ENABLE_MESSAGE_RID_CHECK_ENABLE)
      "TRUE" : TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_BINARY = 1'b1;
      "FALSE" : TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_ENABLE_MESSAGE_RID_CHECK_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", TL_ENABLE_MESSAGE_RID_CHECK_ENABLE);
        #1 $finish;
      end
    endcase

    case (TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE)
      "FALSE" : TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_BINARY = 1'b0;
      "TRUE" : TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE);
        #1 $finish;
      end
    endcase

    case (TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE)
      "FALSE" : TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_BINARY = 1'b0;
      "TRUE" : TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE);
        #1 $finish;
      end
    endcase

    case (TL_LEGACY_MODE_ENABLE)
      "FALSE" : TL_LEGACY_MODE_ENABLE_BINARY = 1'b0;
      "TRUE" : TL_LEGACY_MODE_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_LEGACY_MODE_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_LEGACY_MODE_ENABLE);
        #1 $finish;
      end
    endcase

    case (TL_PF_ENABLE_REG)
      "FALSE" : TL_PF_ENABLE_REG_BINARY = 1'b0;
      "TRUE" : TL_PF_ENABLE_REG_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_PF_ENABLE_REG on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_PF_ENABLE_REG);
        #1 $finish;
      end
    endcase

    case (TL_TAG_MGMT_ENABLE)
      "TRUE" : TL_TAG_MGMT_ENABLE_BINARY = 1'b1;
      "FALSE" : TL_TAG_MGMT_ENABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_TAG_MGMT_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", TL_TAG_MGMT_ENABLE);
        #1 $finish;
      end
    endcase

    case (VF0_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF0_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF0_TPHR_CAP_DEV_SPECIFIC_MODE);
        #1 $finish;
      end
    endcase

    case (VF0_TPHR_CAP_ENABLE)
      "FALSE" : VF0_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF0_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF0_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF0_TPHR_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (VF0_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF0_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF0_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF0_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF0_TPHR_CAP_INT_VEC_MODE);
        #1 $finish;
      end
    endcase

    case (VF1_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF1_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF1_TPHR_CAP_DEV_SPECIFIC_MODE);
        #1 $finish;
      end
    endcase

    case (VF1_TPHR_CAP_ENABLE)
      "FALSE" : VF1_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF1_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF1_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF1_TPHR_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (VF1_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF1_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF1_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF1_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF1_TPHR_CAP_INT_VEC_MODE);
        #1 $finish;
      end
    endcase

    case (VF2_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF2_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF2_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF2_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF2_TPHR_CAP_DEV_SPECIFIC_MODE);
        #1 $finish;
      end
    endcase

    case (VF2_TPHR_CAP_ENABLE)
      "FALSE" : VF2_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF2_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF2_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF2_TPHR_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (VF2_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF2_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF2_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF2_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF2_TPHR_CAP_INT_VEC_MODE);
        #1 $finish;
      end
    endcase

    case (VF3_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF3_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF3_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF3_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF3_TPHR_CAP_DEV_SPECIFIC_MODE);
        #1 $finish;
      end
    endcase

    case (VF3_TPHR_CAP_ENABLE)
      "FALSE" : VF3_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF3_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF3_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF3_TPHR_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (VF3_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF3_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF3_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF3_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF3_TPHR_CAP_INT_VEC_MODE);
        #1 $finish;
      end
    endcase

    case (VF4_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF4_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF4_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF4_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF4_TPHR_CAP_DEV_SPECIFIC_MODE);
        #1 $finish;
      end
    endcase

    case (VF4_TPHR_CAP_ENABLE)
      "FALSE" : VF4_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF4_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF4_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF4_TPHR_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (VF4_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF4_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF4_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF4_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF4_TPHR_CAP_INT_VEC_MODE);
        #1 $finish;
      end
    endcase

    case (VF5_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF5_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF5_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF5_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF5_TPHR_CAP_DEV_SPECIFIC_MODE);
        #1 $finish;
      end
    endcase

    case (VF5_TPHR_CAP_ENABLE)
      "FALSE" : VF5_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF5_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF5_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF5_TPHR_CAP_ENABLE);
        #1 $finish;
      end
    endcase

    case (VF5_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF5_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF5_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF5_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF5_TPHR_CAP_INT_VEC_MODE);
        #1 $finish;
      end
    endcase

    if ((LL_ACK_TIMEOUT_FUNC >= 0) && (LL_ACK_TIMEOUT_FUNC <= 3))
      LL_ACK_TIMEOUT_FUNC_BINARY = LL_ACK_TIMEOUT_FUNC;
    else begin
      $display("Attribute Syntax Error : The Attribute LL_ACK_TIMEOUT_FUNC on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", LL_ACK_TIMEOUT_FUNC);
      #1 $finish;
    end

    if ((LL_REPLAY_TIMEOUT_FUNC >= 0) && (LL_REPLAY_TIMEOUT_FUNC <= 3))
      LL_REPLAY_TIMEOUT_FUNC_BINARY = LL_REPLAY_TIMEOUT_FUNC;
    else begin
      $display("Attribute Syntax Error : The Attribute LL_REPLAY_TIMEOUT_FUNC on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", LL_REPLAY_TIMEOUT_FUNC);
      #1 $finish;
    end

    if ((PF0_DEV_CAP_ENDPOINT_L0S_LATENCY >= 0) && (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY <= 7))
      PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_BINARY = PF0_DEV_CAP_ENDPOINT_L0S_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP_ENDPOINT_L0S_LATENCY on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_DEV_CAP_ENDPOINT_L0S_LATENCY);
      #1 $finish;
    end

    if ((PF0_DEV_CAP_ENDPOINT_L1_LATENCY >= 0) && (PF0_DEV_CAP_ENDPOINT_L1_LATENCY <= 7))
      PF0_DEV_CAP_ENDPOINT_L1_LATENCY_BINARY = PF0_DEV_CAP_ENDPOINT_L1_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP_ENDPOINT_L1_LATENCY on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_DEV_CAP_ENDPOINT_L1_LATENCY);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_ASPM_SUPPORT >= 0) && (PF0_LINK_CAP_ASPM_SUPPORT <= 3))
      PF0_LINK_CAP_ASPM_SUPPORT_BINARY = PF0_LINK_CAP_ASPM_SUPPORT;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_ASPM_SUPPORT on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", PF0_LINK_CAP_ASPM_SUPPORT);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2);
      #1 $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3);
      #1 $finish;
    end

    if ((PF0_MSIX_CAP_PBA_BIR >= 0) && (PF0_MSIX_CAP_PBA_BIR <= 7))
      PF0_MSIX_CAP_PBA_BIR_BINARY = PF0_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_MSIX_CAP_PBA_BIR);
      #1 $finish;
    end

    if ((PF0_MSIX_CAP_TABLE_BIR >= 0) && (PF0_MSIX_CAP_TABLE_BIR <= 7))
      PF0_MSIX_CAP_TABLE_BIR_BINARY = PF0_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_MSIX_CAP_TABLE_BIR);
      #1 $finish;
    end

    if ((PF0_MSI_CAP_MULTIMSGCAP >= 0) && (PF0_MSI_CAP_MULTIMSGCAP <= 7))
      PF0_MSI_CAP_MULTIMSGCAP_BINARY = PF0_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_MSI_CAP_MULTIMSGCAP);
      #1 $finish;
    end

    if ((PF1_MSIX_CAP_PBA_BIR >= 0) && (PF1_MSIX_CAP_PBA_BIR <= 7))
      PF1_MSIX_CAP_PBA_BIR_BINARY = PF1_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute PF1_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF1_MSIX_CAP_PBA_BIR);
      #1 $finish;
    end

    if ((PF1_MSIX_CAP_TABLE_BIR >= 0) && (PF1_MSIX_CAP_TABLE_BIR <= 7))
      PF1_MSIX_CAP_TABLE_BIR_BINARY = PF1_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute PF1_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF1_MSIX_CAP_TABLE_BIR);
      #1 $finish;
    end

    if ((PF1_MSI_CAP_MULTIMSGCAP >= 0) && (PF1_MSI_CAP_MULTIMSGCAP <= 7))
      PF1_MSI_CAP_MULTIMSGCAP_BINARY = PF1_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute PF1_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF1_MSI_CAP_MULTIMSGCAP);
      #1 $finish;
    end

    if ((PL_N_FTS_COMCLK_GEN1 >= 0) && (PL_N_FTS_COMCLK_GEN1 <= 255))
      PL_N_FTS_COMCLK_GEN1_BINARY = PL_N_FTS_COMCLK_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_COMCLK_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_COMCLK_GEN1);
      #1 $finish;
    end

    if ((PL_N_FTS_COMCLK_GEN2 >= 0) && (PL_N_FTS_COMCLK_GEN2 <= 255))
      PL_N_FTS_COMCLK_GEN2_BINARY = PL_N_FTS_COMCLK_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_COMCLK_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_COMCLK_GEN2);
      #1 $finish;
    end

    if ((PL_N_FTS_COMCLK_GEN3 >= 0) && (PL_N_FTS_COMCLK_GEN3 <= 255))
      PL_N_FTS_COMCLK_GEN3_BINARY = PL_N_FTS_COMCLK_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_COMCLK_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_COMCLK_GEN3);
      #1 $finish;
    end

    if ((PL_N_FTS_GEN1 >= 0) && (PL_N_FTS_GEN1 <= 255))
      PL_N_FTS_GEN1_BINARY = PL_N_FTS_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_GEN1);
      #1 $finish;
    end

    if ((PL_N_FTS_GEN2 >= 0) && (PL_N_FTS_GEN2 <= 255))
      PL_N_FTS_GEN2_BINARY = PL_N_FTS_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_GEN2);
      #1 $finish;
    end

    if ((PL_N_FTS_GEN3 >= 0) && (PL_N_FTS_GEN3 <= 255))
      PL_N_FTS_GEN3_BINARY = PL_N_FTS_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_GEN3);
      #1 $finish;
    end

    if ((SPARE_BIT0 >= 0) && (SPARE_BIT0 <= 1))
      SPARE_BIT0_BINARY = SPARE_BIT0;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT0 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT0);
      #1 $finish;
    end

    if ((SPARE_BIT1 >= 0) && (SPARE_BIT1 <= 1))
      SPARE_BIT1_BINARY = SPARE_BIT1;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT1);
      #1 $finish;
    end

    if ((SPARE_BIT2 >= 0) && (SPARE_BIT2 <= 1))
      SPARE_BIT2_BINARY = SPARE_BIT2;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT2);
      #1 $finish;
    end

    if ((SPARE_BIT3 >= 0) && (SPARE_BIT3 <= 1))
      SPARE_BIT3_BINARY = SPARE_BIT3;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT3);
      #1 $finish;
    end

    if ((SPARE_BIT4 >= 0) && (SPARE_BIT4 <= 1))
      SPARE_BIT4_BINARY = SPARE_BIT4;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT4 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT4);
      #1 $finish;
    end

    if ((SPARE_BIT5 >= 0) && (SPARE_BIT5 <= 1))
      SPARE_BIT5_BINARY = SPARE_BIT5;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT5 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT5);
      #1 $finish;
    end

    if ((SPARE_BIT6 >= 0) && (SPARE_BIT6 <= 1))
      SPARE_BIT6_BINARY = SPARE_BIT6;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT6 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT6);
      #1 $finish;
    end

    if ((SPARE_BIT7 >= 0) && (SPARE_BIT7 <= 1))
      SPARE_BIT7_BINARY = SPARE_BIT7;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT7 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT7);
      #1 $finish;
    end

    if ((SPARE_BIT8 >= 0) && (SPARE_BIT8 <= 1))
      SPARE_BIT8_BINARY = SPARE_BIT8;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT8 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT8);
      #1 $finish;
    end

    if ((VF0_MSIX_CAP_PBA_BIR >= 0) && (VF0_MSIX_CAP_PBA_BIR <= 7))
      VF0_MSIX_CAP_PBA_BIR_BINARY = VF0_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF0_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF0_MSIX_CAP_PBA_BIR);
      #1 $finish;
    end

    if ((VF0_MSIX_CAP_TABLE_BIR >= 0) && (VF0_MSIX_CAP_TABLE_BIR <= 7))
      VF0_MSIX_CAP_TABLE_BIR_BINARY = VF0_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF0_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF0_MSIX_CAP_TABLE_BIR);
      #1 $finish;
    end

    if ((VF0_MSI_CAP_MULTIMSGCAP >= 0) && (VF0_MSI_CAP_MULTIMSGCAP <= 7))
      VF0_MSI_CAP_MULTIMSGCAP_BINARY = VF0_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF0_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF0_MSI_CAP_MULTIMSGCAP);
      #1 $finish;
    end

    if ((VF1_MSIX_CAP_PBA_BIR >= 0) && (VF1_MSIX_CAP_PBA_BIR <= 7))
      VF1_MSIX_CAP_PBA_BIR_BINARY = VF1_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF1_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF1_MSIX_CAP_PBA_BIR);
      #1 $finish;
    end

    if ((VF1_MSIX_CAP_TABLE_BIR >= 0) && (VF1_MSIX_CAP_TABLE_BIR <= 7))
      VF1_MSIX_CAP_TABLE_BIR_BINARY = VF1_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF1_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF1_MSIX_CAP_TABLE_BIR);
      #1 $finish;
    end

    if ((VF1_MSI_CAP_MULTIMSGCAP >= 0) && (VF1_MSI_CAP_MULTIMSGCAP <= 7))
      VF1_MSI_CAP_MULTIMSGCAP_BINARY = VF1_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF1_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF1_MSI_CAP_MULTIMSGCAP);
      #1 $finish;
    end

    if ((VF2_MSIX_CAP_PBA_BIR >= 0) && (VF2_MSIX_CAP_PBA_BIR <= 7))
      VF2_MSIX_CAP_PBA_BIR_BINARY = VF2_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF2_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF2_MSIX_CAP_PBA_BIR);
      #1 $finish;
    end

    if ((VF2_MSIX_CAP_TABLE_BIR >= 0) && (VF2_MSIX_CAP_TABLE_BIR <= 7))
      VF2_MSIX_CAP_TABLE_BIR_BINARY = VF2_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF2_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF2_MSIX_CAP_TABLE_BIR);
      #1 $finish;
    end

    if ((VF2_MSI_CAP_MULTIMSGCAP >= 0) && (VF2_MSI_CAP_MULTIMSGCAP <= 7))
      VF2_MSI_CAP_MULTIMSGCAP_BINARY = VF2_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF2_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF2_MSI_CAP_MULTIMSGCAP);
      #1 $finish;
    end

    if ((VF3_MSIX_CAP_PBA_BIR >= 0) && (VF3_MSIX_CAP_PBA_BIR <= 7))
      VF3_MSIX_CAP_PBA_BIR_BINARY = VF3_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF3_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF3_MSIX_CAP_PBA_BIR);
      #1 $finish;
    end

    if ((VF3_MSIX_CAP_TABLE_BIR >= 0) && (VF3_MSIX_CAP_TABLE_BIR <= 7))
      VF3_MSIX_CAP_TABLE_BIR_BINARY = VF3_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF3_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF3_MSIX_CAP_TABLE_BIR);
      #1 $finish;
    end

    if ((VF3_MSI_CAP_MULTIMSGCAP >= 0) && (VF3_MSI_CAP_MULTIMSGCAP <= 7))
      VF3_MSI_CAP_MULTIMSGCAP_BINARY = VF3_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF3_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF3_MSI_CAP_MULTIMSGCAP);
      #1 $finish;
    end

    if ((VF4_MSIX_CAP_PBA_BIR >= 0) && (VF4_MSIX_CAP_PBA_BIR <= 7))
      VF4_MSIX_CAP_PBA_BIR_BINARY = VF4_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF4_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF4_MSIX_CAP_PBA_BIR);
      #1 $finish;
    end

    if ((VF4_MSIX_CAP_TABLE_BIR >= 0) && (VF4_MSIX_CAP_TABLE_BIR <= 7))
      VF4_MSIX_CAP_TABLE_BIR_BINARY = VF4_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF4_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF4_MSIX_CAP_TABLE_BIR);
      #1 $finish;
    end

    if ((VF4_MSI_CAP_MULTIMSGCAP >= 0) && (VF4_MSI_CAP_MULTIMSGCAP <= 7))
      VF4_MSI_CAP_MULTIMSGCAP_BINARY = VF4_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF4_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF4_MSI_CAP_MULTIMSGCAP);
      #1 $finish;
    end

    if ((VF5_MSIX_CAP_PBA_BIR >= 0) && (VF5_MSIX_CAP_PBA_BIR <= 7))
      VF5_MSIX_CAP_PBA_BIR_BINARY = VF5_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF5_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF5_MSIX_CAP_PBA_BIR);
      #1 $finish;
    end

    if ((VF5_MSIX_CAP_TABLE_BIR >= 0) && (VF5_MSIX_CAP_TABLE_BIR <= 7))
      VF5_MSIX_CAP_TABLE_BIR_BINARY = VF5_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF5_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF5_MSIX_CAP_TABLE_BIR);
      #1 $finish;
    end

    if ((VF5_MSI_CAP_MULTIMSGCAP >= 0) && (VF5_MSI_CAP_MULTIMSGCAP <= 7))
      VF5_MSI_CAP_MULTIMSGCAP_BINARY = VF5_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF5_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF5_MSI_CAP_MULTIMSGCAP);
      #1 $finish;
    end

  end

  wire [11:0] delay_CFGFCCPLD;
  wire [11:0] delay_CFGFCNPD;
  wire [11:0] delay_CFGFCPD;
  wire [11:0] delay_CFGVFSTATUS;
  wire [143:0] delay_MIREPLAYRAMWRITEDATA;
  wire [143:0] delay_MIREQUESTRAMWRITEDATA;
  wire [15:0] delay_CFGPERFUNCSTATUSDATA;
  wire [15:0] delay_DBGDATAOUT;
  wire [15:0] delay_DRPDO;
  wire [17:0] delay_CFGVFPOWERSTATE;
  wire [17:0] delay_CFGVFTPHSTMODE;
  wire [1:0] delay_CFGDPASUBSTATECHANGE;
  wire [1:0] delay_CFGFLRINPROCESS;
  wire [1:0] delay_CFGINTERRUPTMSIENABLE;
  wire [1:0] delay_CFGINTERRUPTMSIXENABLE;
  wire [1:0] delay_CFGINTERRUPTMSIXMASK;
  wire [1:0] delay_CFGLINKPOWERSTATE;
  wire [1:0] delay_CFGOBFFENABLE;
  wire [1:0] delay_CFGPHYLINKSTATUS;
  wire [1:0] delay_CFGRCBSTATUS;
  wire [1:0] delay_CFGTPHREQUESTERENABLE;
  wire [1:0] delay_MIREPLAYRAMREADENABLE;
  wire [1:0] delay_MIREPLAYRAMWRITEENABLE;
  wire [1:0] delay_PCIERQTAGAV;
  wire [1:0] delay_PCIETFCNPDAV;
  wire [1:0] delay_PCIETFCNPHAV;
  wire [1:0] delay_PIPERX0EQCONTROL;
  wire [1:0] delay_PIPERX1EQCONTROL;
  wire [1:0] delay_PIPERX2EQCONTROL;
  wire [1:0] delay_PIPERX3EQCONTROL;
  wire [1:0] delay_PIPERX4EQCONTROL;
  wire [1:0] delay_PIPERX5EQCONTROL;
  wire [1:0] delay_PIPERX6EQCONTROL;
  wire [1:0] delay_PIPERX7EQCONTROL;
  wire [1:0] delay_PIPETX0CHARISK;
  wire [1:0] delay_PIPETX0EQCONTROL;
  wire [1:0] delay_PIPETX0POWERDOWN;
  wire [1:0] delay_PIPETX0SYNCHEADER;
  wire [1:0] delay_PIPETX1CHARISK;
  wire [1:0] delay_PIPETX1EQCONTROL;
  wire [1:0] delay_PIPETX1POWERDOWN;
  wire [1:0] delay_PIPETX1SYNCHEADER;
  wire [1:0] delay_PIPETX2CHARISK;
  wire [1:0] delay_PIPETX2EQCONTROL;
  wire [1:0] delay_PIPETX2POWERDOWN;
  wire [1:0] delay_PIPETX2SYNCHEADER;
  wire [1:0] delay_PIPETX3CHARISK;
  wire [1:0] delay_PIPETX3EQCONTROL;
  wire [1:0] delay_PIPETX3POWERDOWN;
  wire [1:0] delay_PIPETX3SYNCHEADER;
  wire [1:0] delay_PIPETX4CHARISK;
  wire [1:0] delay_PIPETX4EQCONTROL;
  wire [1:0] delay_PIPETX4POWERDOWN;
  wire [1:0] delay_PIPETX4SYNCHEADER;
  wire [1:0] delay_PIPETX5CHARISK;
  wire [1:0] delay_PIPETX5EQCONTROL;
  wire [1:0] delay_PIPETX5POWERDOWN;
  wire [1:0] delay_PIPETX5SYNCHEADER;
  wire [1:0] delay_PIPETX6CHARISK;
  wire [1:0] delay_PIPETX6EQCONTROL;
  wire [1:0] delay_PIPETX6POWERDOWN;
  wire [1:0] delay_PIPETX6SYNCHEADER;
  wire [1:0] delay_PIPETX7CHARISK;
  wire [1:0] delay_PIPETX7EQCONTROL;
  wire [1:0] delay_PIPETX7POWERDOWN;
  wire [1:0] delay_PIPETX7SYNCHEADER;
  wire [1:0] delay_PIPETXRATE;
  wire [1:0] delay_PLEQPHASE;
  wire [255:0] delay_MAXISCQTDATA;
  wire [255:0] delay_MAXISRCTDATA;
  wire [2:0] delay_CFGCURRENTSPEED;
  wire [2:0] delay_CFGMAXPAYLOAD;
  wire [2:0] delay_CFGMAXREADREQ;
  wire [2:0] delay_CFGTPHFUNCTIONNUM;
  wire [2:0] delay_PIPERX0EQPRESET;
  wire [2:0] delay_PIPERX1EQPRESET;
  wire [2:0] delay_PIPERX2EQPRESET;
  wire [2:0] delay_PIPERX3EQPRESET;
  wire [2:0] delay_PIPERX4EQPRESET;
  wire [2:0] delay_PIPERX5EQPRESET;
  wire [2:0] delay_PIPERX6EQPRESET;
  wire [2:0] delay_PIPERX7EQPRESET;
  wire [2:0] delay_PIPETXMARGIN;
  wire [31:0] delay_CFGEXTWRITEDATA;
  wire [31:0] delay_CFGINTERRUPTMSIDATA;
  wire [31:0] delay_CFGMGMTREADDATA;
  wire [31:0] delay_CFGTPHSTTWRITEDATA;
  wire [31:0] delay_PIPETX0DATA;
  wire [31:0] delay_PIPETX1DATA;
  wire [31:0] delay_PIPETX2DATA;
  wire [31:0] delay_PIPETX3DATA;
  wire [31:0] delay_PIPETX4DATA;
  wire [31:0] delay_PIPETX5DATA;
  wire [31:0] delay_PIPETX6DATA;
  wire [31:0] delay_PIPETX7DATA;
  wire [3:0] delay_CFGEXTWRITEBYTEENABLE;
  wire [3:0] delay_CFGNEGOTIATEDWIDTH;
  wire [3:0] delay_CFGTPHSTTWRITEBYTEVALID;
  wire [3:0] delay_MICOMPLETIONRAMREADENABLEL;
  wire [3:0] delay_MICOMPLETIONRAMREADENABLEU;
  wire [3:0] delay_MICOMPLETIONRAMWRITEENABLEL;
  wire [3:0] delay_MICOMPLETIONRAMWRITEENABLEU;
  wire [3:0] delay_MIREQUESTRAMREADENABLE;
  wire [3:0] delay_MIREQUESTRAMWRITEENABLE;
  wire [3:0] delay_PCIERQSEQNUM;
  wire [3:0] delay_PIPERX0EQLPTXPRESET;
  wire [3:0] delay_PIPERX1EQLPTXPRESET;
  wire [3:0] delay_PIPERX2EQLPTXPRESET;
  wire [3:0] delay_PIPERX3EQLPTXPRESET;
  wire [3:0] delay_PIPERX4EQLPTXPRESET;
  wire [3:0] delay_PIPERX5EQLPTXPRESET;
  wire [3:0] delay_PIPERX6EQLPTXPRESET;
  wire [3:0] delay_PIPERX7EQLPTXPRESET;
  wire [3:0] delay_PIPETX0EQPRESET;
  wire [3:0] delay_PIPETX1EQPRESET;
  wire [3:0] delay_PIPETX2EQPRESET;
  wire [3:0] delay_PIPETX3EQPRESET;
  wire [3:0] delay_PIPETX4EQPRESET;
  wire [3:0] delay_PIPETX5EQPRESET;
  wire [3:0] delay_PIPETX6EQPRESET;
  wire [3:0] delay_PIPETX7EQPRESET;
  wire [3:0] delay_SAXISCCTREADY;
  wire [3:0] delay_SAXISRQTREADY;
  wire [4:0] delay_CFGMSGRECEIVEDTYPE;
  wire [4:0] delay_CFGTPHSTTADDRESS;
  wire [5:0] delay_CFGFUNCTIONPOWERSTATE;
  wire [5:0] delay_CFGINTERRUPTMSIMMENABLE;
  wire [5:0] delay_CFGINTERRUPTMSIVFENABLE;
  wire [5:0] delay_CFGINTERRUPTMSIXVFENABLE;
  wire [5:0] delay_CFGINTERRUPTMSIXVFMASK;
  wire [5:0] delay_CFGLTSSMSTATE;
  wire [5:0] delay_CFGTPHSTMODE;
  wire [5:0] delay_CFGVFFLRINPROCESS;
  wire [5:0] delay_CFGVFTPHREQUESTERENABLE;
  wire [5:0] delay_PCIECQNPREQCOUNT;
  wire [5:0] delay_PCIERQTAG;
  wire [5:0] delay_PIPERX0EQLPLFFS;
  wire [5:0] delay_PIPERX1EQLPLFFS;
  wire [5:0] delay_PIPERX2EQLPLFFS;
  wire [5:0] delay_PIPERX3EQLPLFFS;
  wire [5:0] delay_PIPERX4EQLPLFFS;
  wire [5:0] delay_PIPERX5EQLPLFFS;
  wire [5:0] delay_PIPERX6EQLPLFFS;
  wire [5:0] delay_PIPERX7EQLPLFFS;
  wire [5:0] delay_PIPETX0EQDEEMPH;
  wire [5:0] delay_PIPETX1EQDEEMPH;
  wire [5:0] delay_PIPETX2EQDEEMPH;
  wire [5:0] delay_PIPETX3EQDEEMPH;
  wire [5:0] delay_PIPETX4EQDEEMPH;
  wire [5:0] delay_PIPETX5EQDEEMPH;
  wire [5:0] delay_PIPETX6EQDEEMPH;
  wire [5:0] delay_PIPETX7EQDEEMPH;
  wire [71:0] delay_MICOMPLETIONRAMWRITEDATAL;
  wire [71:0] delay_MICOMPLETIONRAMWRITEDATAU;
  wire [74:0] delay_MAXISRCTUSER;
  wire [7:0] delay_CFGEXTFUNCTIONNUMBER;
  wire [7:0] delay_CFGFCCPLH;
  wire [7:0] delay_CFGFCNPH;
  wire [7:0] delay_CFGFCPH;
  wire [7:0] delay_CFGFUNCTIONSTATUS;
  wire [7:0] delay_CFGMSGRECEIVEDDATA;
  wire [7:0] delay_MAXISCQTKEEP;
  wire [7:0] delay_MAXISRCTKEEP;
  wire [7:0] delay_PLGEN3PCSRXSLIDE;
  wire [84:0] delay_MAXISCQTUSER;
  wire [8:0] delay_MIREPLAYRAMADDRESS;
  wire [8:0] delay_MIREQUESTRAMREADADDRESSA;
  wire [8:0] delay_MIREQUESTRAMREADADDRESSB;
  wire [8:0] delay_MIREQUESTRAMWRITEADDRESSA;
  wire [8:0] delay_MIREQUESTRAMWRITEADDRESSB;
  wire [9:0] delay_CFGEXTREGISTERNUMBER;
  wire [9:0] delay_MICOMPLETIONRAMREADADDRESSAL;
  wire [9:0] delay_MICOMPLETIONRAMREADADDRESSAU;
  wire [9:0] delay_MICOMPLETIONRAMREADADDRESSBL;
  wire [9:0] delay_MICOMPLETIONRAMREADADDRESSBU;
  wire [9:0] delay_MICOMPLETIONRAMWRITEADDRESSAL;
  wire [9:0] delay_MICOMPLETIONRAMWRITEADDRESSAU;
  wire [9:0] delay_MICOMPLETIONRAMWRITEADDRESSBL;
  wire [9:0] delay_MICOMPLETIONRAMWRITEADDRESSBU;
  wire delay_CFGERRCOROUT;
  wire delay_CFGERRFATALOUT;
  wire delay_CFGERRNONFATALOUT;
  wire delay_CFGEXTREADRECEIVED;
  wire delay_CFGEXTWRITERECEIVED;
  wire delay_CFGHOTRESETOUT;
  wire delay_CFGINPUTUPDATEDONE;
  wire delay_CFGINTERRUPTAOUTPUT;
  wire delay_CFGINTERRUPTBOUTPUT;
  wire delay_CFGINTERRUPTCOUTPUT;
  wire delay_CFGINTERRUPTDOUTPUT;
  wire delay_CFGINTERRUPTMSIFAIL;
  wire delay_CFGINTERRUPTMSIMASKUPDATE;
  wire delay_CFGINTERRUPTMSISENT;
  wire delay_CFGINTERRUPTMSIXFAIL;
  wire delay_CFGINTERRUPTMSIXSENT;
  wire delay_CFGINTERRUPTSENT;
  wire delay_CFGLOCALERROR;
  wire delay_CFGLTRENABLE;
  wire delay_CFGMCUPDATEDONE;
  wire delay_CFGMGMTREADWRITEDONE;
  wire delay_CFGMSGRECEIVED;
  wire delay_CFGMSGTRANSMITDONE;
  wire delay_CFGPERFUNCTIONUPDATEDONE;
  wire delay_CFGPHYLINKDOWN;
  wire delay_CFGPLSTATUSCHANGE;
  wire delay_CFGPOWERSTATECHANGEINTERRUPT;
  wire delay_CFGTPHSTTREADENABLE;
  wire delay_CFGTPHSTTWRITEENABLE;
  wire delay_DRPRDY;
  wire delay_MAXISCQTLAST;
  wire delay_MAXISCQTVALID;
  wire delay_MAXISRCTLAST;
  wire delay_MAXISRCTVALID;
  wire delay_PCIERQSEQNUMVLD;
  wire delay_PCIERQTAGVLD;
  wire delay_PIPERX0POLARITY;
  wire delay_PIPERX1POLARITY;
  wire delay_PIPERX2POLARITY;
  wire delay_PIPERX3POLARITY;
  wire delay_PIPERX4POLARITY;
  wire delay_PIPERX5POLARITY;
  wire delay_PIPERX6POLARITY;
  wire delay_PIPERX7POLARITY;
  wire delay_PIPETX0COMPLIANCE;
  wire delay_PIPETX0DATAVALID;
  wire delay_PIPETX0ELECIDLE;
  wire delay_PIPETX0STARTBLOCK;
  wire delay_PIPETX1COMPLIANCE;
  wire delay_PIPETX1DATAVALID;
  wire delay_PIPETX1ELECIDLE;
  wire delay_PIPETX1STARTBLOCK;
  wire delay_PIPETX2COMPLIANCE;
  wire delay_PIPETX2DATAVALID;
  wire delay_PIPETX2ELECIDLE;
  wire delay_PIPETX2STARTBLOCK;
  wire delay_PIPETX3COMPLIANCE;
  wire delay_PIPETX3DATAVALID;
  wire delay_PIPETX3ELECIDLE;
  wire delay_PIPETX3STARTBLOCK;
  wire delay_PIPETX4COMPLIANCE;
  wire delay_PIPETX4DATAVALID;
  wire delay_PIPETX4ELECIDLE;
  wire delay_PIPETX4STARTBLOCK;
  wire delay_PIPETX5COMPLIANCE;
  wire delay_PIPETX5DATAVALID;
  wire delay_PIPETX5ELECIDLE;
  wire delay_PIPETX5STARTBLOCK;
  wire delay_PIPETX6COMPLIANCE;
  wire delay_PIPETX6DATAVALID;
  wire delay_PIPETX6ELECIDLE;
  wire delay_PIPETX6STARTBLOCK;
  wire delay_PIPETX7COMPLIANCE;
  wire delay_PIPETX7DATAVALID;
  wire delay_PIPETX7ELECIDLE;
  wire delay_PIPETX7STARTBLOCK;
  wire delay_PIPETXDEEMPH;
  wire delay_PIPETXRCVRDET;
  wire delay_PIPETXRESET;
  wire delay_PIPETXSWING;
  wire delay_PLEQINPROGRESS;

  wire [10:0] delay_DRPADDR;
  wire [143:0] delay_MICOMPLETIONRAMREADDATA;
  wire [143:0] delay_MIREPLAYRAMREADDATA;
  wire [143:0] delay_MIREQUESTRAMREADDATA;
  wire [15:0] delay_CFGDEVID;
  wire [15:0] delay_CFGSUBSYSID;
  wire [15:0] delay_CFGSUBSYSVENDID;
  wire [15:0] delay_CFGVENDID;
  wire [15:0] delay_DRPDI;
  wire [17:0] delay_PIPERX0EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX1EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX2EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX3EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX4EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX5EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX6EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX7EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPETX0EQCOEFF;
  wire [17:0] delay_PIPETX1EQCOEFF;
  wire [17:0] delay_PIPETX2EQCOEFF;
  wire [17:0] delay_PIPETX3EQCOEFF;
  wire [17:0] delay_PIPETX4EQCOEFF;
  wire [17:0] delay_PIPETX5EQCOEFF;
  wire [17:0] delay_PIPETX6EQCOEFF;
  wire [17:0] delay_PIPETX7EQCOEFF;
  wire [18:0] delay_CFGMGMTADDR;
  wire [1:0] delay_CFGFLRDONE;
  wire [1:0] delay_CFGINTERRUPTMSITPHTYPE;
  wire [1:0] delay_CFGINTERRUPTPENDING;
  wire [1:0] delay_PIPERX0CHARISK;
  wire [1:0] delay_PIPERX0SYNCHEADER;
  wire [1:0] delay_PIPERX1CHARISK;
  wire [1:0] delay_PIPERX1SYNCHEADER;
  wire [1:0] delay_PIPERX2CHARISK;
  wire [1:0] delay_PIPERX2SYNCHEADER;
  wire [1:0] delay_PIPERX3CHARISK;
  wire [1:0] delay_PIPERX3SYNCHEADER;
  wire [1:0] delay_PIPERX4CHARISK;
  wire [1:0] delay_PIPERX4SYNCHEADER;
  wire [1:0] delay_PIPERX5CHARISK;
  wire [1:0] delay_PIPERX5SYNCHEADER;
  wire [1:0] delay_PIPERX6CHARISK;
  wire [1:0] delay_PIPERX6SYNCHEADER;
  wire [1:0] delay_PIPERX7CHARISK;
  wire [1:0] delay_PIPERX7SYNCHEADER;
  wire [21:0] delay_MAXISCQTREADY;
  wire [21:0] delay_MAXISRCTREADY;
  wire [255:0] delay_SAXISCCTDATA;
  wire [255:0] delay_SAXISRQTDATA;
  wire [2:0] delay_CFGDSFUNCTIONNUMBER;
  wire [2:0] delay_CFGFCSEL;
  wire [2:0] delay_CFGINTERRUPTMSIATTR;
  wire [2:0] delay_CFGINTERRUPTMSIFUNCTIONNUMBER;
  wire [2:0] delay_CFGMSGTRANSMITTYPE;
  wire [2:0] delay_CFGPERFUNCSTATUSCONTROL;
  wire [2:0] delay_CFGPERFUNCTIONNUMBER;
  wire [2:0] delay_PIPERX0STATUS;
  wire [2:0] delay_PIPERX1STATUS;
  wire [2:0] delay_PIPERX2STATUS;
  wire [2:0] delay_PIPERX3STATUS;
  wire [2:0] delay_PIPERX4STATUS;
  wire [2:0] delay_PIPERX5STATUS;
  wire [2:0] delay_PIPERX6STATUS;
  wire [2:0] delay_PIPERX7STATUS;
  wire [31:0] delay_CFGEXTREADDATA;
  wire [31:0] delay_CFGINTERRUPTMSIINT;
  wire [31:0] delay_CFGINTERRUPTMSIXDATA;
  wire [31:0] delay_CFGMGMTWRITEDATA;
  wire [31:0] delay_CFGMSGTRANSMITDATA;
  wire [31:0] delay_CFGTPHSTTREADDATA;
  wire [31:0] delay_PIPERX0DATA;
  wire [31:0] delay_PIPERX1DATA;
  wire [31:0] delay_PIPERX2DATA;
  wire [31:0] delay_PIPERX3DATA;
  wire [31:0] delay_PIPERX4DATA;
  wire [31:0] delay_PIPERX5DATA;
  wire [31:0] delay_PIPERX6DATA;
  wire [31:0] delay_PIPERX7DATA;
  wire [32:0] delay_SAXISCCTUSER;
  wire [3:0] delay_CFGINTERRUPTINT;
  wire [3:0] delay_CFGINTERRUPTMSISELECT;
  wire [3:0] delay_CFGMGMTBYTEENABLE;
  wire [4:0] delay_CFGDSDEVICENUMBER;
  wire [59:0] delay_SAXISRQTUSER;
  wire [5:0] delay_CFGVFFLRDONE;
  wire [5:0] delay_PIPEEQFS;
  wire [5:0] delay_PIPEEQLF;
  wire [63:0] delay_CFGDSN;
  wire [63:0] delay_CFGINTERRUPTMSIPENDINGSTATUS;
  wire [63:0] delay_CFGINTERRUPTMSIXADDRESS;
  wire [7:0] delay_CFGDSBUSNUMBER;
  wire [7:0] delay_CFGDSPORTNUMBER;
  wire [7:0] delay_CFGREVID;
  wire [7:0] delay_PLGEN3PCSRXSYNCDONE;
  wire [7:0] delay_SAXISCCTKEEP;
  wire [7:0] delay_SAXISRQTKEEP;
  wire [8:0] delay_CFGINTERRUPTMSITPHSTTAG;
  wire delay_CFGCONFIGSPACEENABLE;
  wire delay_CFGERRCORIN;
  wire delay_CFGERRUNCORIN;
  wire delay_CFGEXTREADDATAVALID;
  wire delay_CFGHOTRESETIN;
  wire delay_CFGINPUTUPDATEREQUEST;
  wire delay_CFGINTERRUPTMSITPHPRESENT;
  wire delay_CFGINTERRUPTMSIXINT;
  wire delay_CFGLINKTRAININGENABLE;
  wire delay_CFGMCUPDATEREQUEST;
  wire delay_CFGMGMTREAD;
  wire delay_CFGMGMTTYPE1CFGREGACCESS;
  wire delay_CFGMGMTWRITE;
  wire delay_CFGMSGTRANSMIT;
  wire delay_CFGPERFUNCTIONOUTPUTREQUEST;
  wire delay_CFGPOWERSTATECHANGEACK;
  wire delay_CFGREQPMTRANSITIONL23READY;
  wire delay_CFGTPHSTTREADDATAVALID;
  wire delay_CORECLK;
  wire delay_CORECLKMICOMPLETIONRAML;
  wire delay_CORECLKMICOMPLETIONRAMU;
  wire delay_CORECLKMIREPLAYRAM;
  wire delay_CORECLKMIREQUESTRAM;
  wire delay_DRPCLK;
  wire delay_DRPEN;
  wire delay_DRPWE;
  wire delay_MGMTRESETN;
  wire delay_MGMTSTICKYRESETN;
  wire delay_PCIECQNPREQ;
  wire delay_PIPECLK;
  wire delay_PIPERESETN;
  wire delay_PIPERX0DATAVALID;
  wire delay_PIPERX0ELECIDLE;
  wire delay_PIPERX0EQDONE;
  wire delay_PIPERX0EQLPADAPTDONE;
  wire delay_PIPERX0EQLPLFFSSEL;
  wire delay_PIPERX0PHYSTATUS;
  wire delay_PIPERX0STARTBLOCK;
  wire delay_PIPERX0VALID;
  wire delay_PIPERX1DATAVALID;
  wire delay_PIPERX1ELECIDLE;
  wire delay_PIPERX1EQDONE;
  wire delay_PIPERX1EQLPADAPTDONE;
  wire delay_PIPERX1EQLPLFFSSEL;
  wire delay_PIPERX1PHYSTATUS;
  wire delay_PIPERX1STARTBLOCK;
  wire delay_PIPERX1VALID;
  wire delay_PIPERX2DATAVALID;
  wire delay_PIPERX2ELECIDLE;
  wire delay_PIPERX2EQDONE;
  wire delay_PIPERX2EQLPADAPTDONE;
  wire delay_PIPERX2EQLPLFFSSEL;
  wire delay_PIPERX2PHYSTATUS;
  wire delay_PIPERX2STARTBLOCK;
  wire delay_PIPERX2VALID;
  wire delay_PIPERX3DATAVALID;
  wire delay_PIPERX3ELECIDLE;
  wire delay_PIPERX3EQDONE;
  wire delay_PIPERX3EQLPADAPTDONE;
  wire delay_PIPERX3EQLPLFFSSEL;
  wire delay_PIPERX3PHYSTATUS;
  wire delay_PIPERX3STARTBLOCK;
  wire delay_PIPERX3VALID;
  wire delay_PIPERX4DATAVALID;
  wire delay_PIPERX4ELECIDLE;
  wire delay_PIPERX4EQDONE;
  wire delay_PIPERX4EQLPADAPTDONE;
  wire delay_PIPERX4EQLPLFFSSEL;
  wire delay_PIPERX4PHYSTATUS;
  wire delay_PIPERX4STARTBLOCK;
  wire delay_PIPERX4VALID;
  wire delay_PIPERX5DATAVALID;
  wire delay_PIPERX5ELECIDLE;
  wire delay_PIPERX5EQDONE;
  wire delay_PIPERX5EQLPADAPTDONE;
  wire delay_PIPERX5EQLPLFFSSEL;
  wire delay_PIPERX5PHYSTATUS;
  wire delay_PIPERX5STARTBLOCK;
  wire delay_PIPERX5VALID;
  wire delay_PIPERX6DATAVALID;
  wire delay_PIPERX6ELECIDLE;
  wire delay_PIPERX6EQDONE;
  wire delay_PIPERX6EQLPADAPTDONE;
  wire delay_PIPERX6EQLPLFFSSEL;
  wire delay_PIPERX6PHYSTATUS;
  wire delay_PIPERX6STARTBLOCK;
  wire delay_PIPERX6VALID;
  wire delay_PIPERX7DATAVALID;
  wire delay_PIPERX7ELECIDLE;
  wire delay_PIPERX7EQDONE;
  wire delay_PIPERX7EQLPADAPTDONE;
  wire delay_PIPERX7EQLPLFFSSEL;
  wire delay_PIPERX7PHYSTATUS;
  wire delay_PIPERX7STARTBLOCK;
  wire delay_PIPERX7VALID;
  wire delay_PIPETX0EQDONE;
  wire delay_PIPETX1EQDONE;
  wire delay_PIPETX2EQDONE;
  wire delay_PIPETX3EQDONE;
  wire delay_PIPETX4EQDONE;
  wire delay_PIPETX5EQDONE;
  wire delay_PIPETX6EQDONE;
  wire delay_PIPETX7EQDONE;
  wire delay_PLDISABLESCRAMBLER;
  wire delay_PLEQRESETEIEOSCOUNT;
  wire delay_PLGEN3PCSDISABLE;
  wire delay_RECCLK;
  wire delay_RESETN;
  wire delay_SAXISCCTLAST;
  wire delay_SAXISCCTVALID;
  wire delay_SAXISRQTLAST;
  wire delay_SAXISRQTVALID;
  wire delay_USERCLK;

   
   //drp monitor
   reg drpen_r1 = 1'b0;
   reg drpen_r2 = 1'b0;
   reg drpwe_r1 = 1'b0;
   reg drpwe_r2 = 1'b0;
   
   reg [1:0] sfsm = 2'b01;
    
   localparam FSM_IDLE = 2'b01;  
   localparam FSM_WAIT = 2'b10;
  

   always @(posedge delay_DRPCLK)
     begin
	// pipeline the DRPEN and DRPWE
        drpen_r1 <= delay_DRPEN;
        drpwe_r1 <= delay_DRPWE;
	drpen_r2 <= drpen_r1;
        drpwe_r2 <= drpwe_r1;

	
	// Check -  if DRPEN or DRPWE is more than 1 DCLK
	if ((drpen_r1 == 1'b1) && (drpen_r2 == 1'b1)) 
	  begin
	     $display("DRC Error : DRPEN is high for more than 1 DRPCLK on %m instance");
	     $finish; 
          end
	
	if ((drpwe_r1 == 1'b1) && (drpwe_r2 == 1'b1))
	  begin
             $display("DRC Error : DRPWE is high for more than 1 DRPCLK on %m instance");
             $finish;
          end


	//After the 1st DRPEN pulse, check the DRPEN and DRPRDY.
	case (sfsm)
          FSM_IDLE:   
            begin
               if(delay_DRPEN == 1'b1)
		 sfsm <= FSM_WAIT;  
            end
          
          FSM_WAIT:
            begin
               // After the 1st DRPEN, 4 cases can happen
               // DRPEN DRPRDY NEXT STATE
               // 0     0      FSM_WAIT - wait for DRPRDY
               // 0     1      FSM_IDLE - normal operation
               // 1     0      FSM_WAIT - display error and wait for DRPRDY
               // 1     1      FSM_WAIT - normal operation. Per UG470, DRPEN and DRPRDY can be at the same cycle.
               
               //Add the check for another DPREN pulse
               if(delay_DRPEN === 1'b1 && delay_DRPRDY === 1'b0) 
		 begin
		    $display("DRC Error : DRPEN is enabled before DRPRDY returns on %m instance");  
		    $finish;
		 end

               //Add the check for another DRPWE pulse
               if ((delay_DRPWE === 1'b1) && (delay_DRPEN === 1'b0))
		 begin
		    $display("DRC Error : DRPWE is enabled before DRPRDY returns on %m instance");
		    $finish;
		 end
                    
               if ((delay_DRPRDY === 1'b1) && (delay_DRPEN === 1'b0))
		 begin
		    sfsm <= FSM_IDLE;
		 end  
               
               if ((delay_DRPRDY === 1'b1)&& (delay_DRPEN === 1'b1))
		 begin
		    sfsm <= FSM_WAIT;
		 end  
            end
        
          default:                  
            begin
               $display("DRC Error : Default state in DRP FSM.");
               $finish;
            end
	endcase

     end // always @ (posedge delay_DRPCLK)
   //end drp monitor   

   
  assign #(out_delay) CFGCURRENTSPEED = delay_CFGCURRENTSPEED;
  assign #(out_delay) CFGDPASUBSTATECHANGE = delay_CFGDPASUBSTATECHANGE;
  assign #(out_delay) CFGERRCOROUT = delay_CFGERRCOROUT;
  assign #(out_delay) CFGERRFATALOUT = delay_CFGERRFATALOUT;
  assign #(out_delay) CFGERRNONFATALOUT = delay_CFGERRNONFATALOUT;
  assign #(out_delay) CFGEXTFUNCTIONNUMBER = delay_CFGEXTFUNCTIONNUMBER;
  assign #(out_delay) CFGEXTREADRECEIVED = delay_CFGEXTREADRECEIVED;
  assign #(out_delay) CFGEXTREGISTERNUMBER = delay_CFGEXTREGISTERNUMBER;
  assign #(out_delay) CFGEXTWRITEBYTEENABLE = delay_CFGEXTWRITEBYTEENABLE;
  assign #(out_delay) CFGEXTWRITEDATA = delay_CFGEXTWRITEDATA;
  assign #(out_delay) CFGEXTWRITERECEIVED = delay_CFGEXTWRITERECEIVED;
  assign #(out_delay) CFGFCCPLD = delay_CFGFCCPLD;
  assign #(out_delay) CFGFCCPLH = delay_CFGFCCPLH;
  assign #(out_delay) CFGFCNPD = delay_CFGFCNPD;
  assign #(out_delay) CFGFCNPH = delay_CFGFCNPH;
  assign #(out_delay) CFGFCPD = delay_CFGFCPD;
  assign #(out_delay) CFGFCPH = delay_CFGFCPH;
  assign #(out_delay) CFGFLRINPROCESS = delay_CFGFLRINPROCESS;
  assign #(out_delay) CFGFUNCTIONPOWERSTATE = delay_CFGFUNCTIONPOWERSTATE;
  assign #(out_delay) CFGFUNCTIONSTATUS = delay_CFGFUNCTIONSTATUS;
  assign #(out_delay) CFGHOTRESETOUT = delay_CFGHOTRESETOUT;
  assign #(out_delay) CFGINPUTUPDATEDONE = delay_CFGINPUTUPDATEDONE;
  assign #(out_delay) CFGINTERRUPTAOUTPUT = delay_CFGINTERRUPTAOUTPUT;
  assign #(out_delay) CFGINTERRUPTBOUTPUT = delay_CFGINTERRUPTBOUTPUT;
  assign #(out_delay) CFGINTERRUPTCOUTPUT = delay_CFGINTERRUPTCOUTPUT;
  assign #(out_delay) CFGINTERRUPTDOUTPUT = delay_CFGINTERRUPTDOUTPUT;
  assign #(out_delay) CFGINTERRUPTMSIDATA = delay_CFGINTERRUPTMSIDATA;
  assign #(out_delay) CFGINTERRUPTMSIENABLE = delay_CFGINTERRUPTMSIENABLE;
  assign #(out_delay) CFGINTERRUPTMSIFAIL = delay_CFGINTERRUPTMSIFAIL;
  assign #(out_delay) CFGINTERRUPTMSIMASKUPDATE = delay_CFGINTERRUPTMSIMASKUPDATE;
  assign #(out_delay) CFGINTERRUPTMSIMMENABLE = delay_CFGINTERRUPTMSIMMENABLE;
  assign #(out_delay) CFGINTERRUPTMSISENT = delay_CFGINTERRUPTMSISENT;
  assign #(out_delay) CFGINTERRUPTMSIVFENABLE = delay_CFGINTERRUPTMSIVFENABLE;
  assign #(out_delay) CFGINTERRUPTMSIXENABLE = delay_CFGINTERRUPTMSIXENABLE;
  assign #(out_delay) CFGINTERRUPTMSIXFAIL = delay_CFGINTERRUPTMSIXFAIL;
  assign #(out_delay) CFGINTERRUPTMSIXMASK = delay_CFGINTERRUPTMSIXMASK;
  assign #(out_delay) CFGINTERRUPTMSIXSENT = delay_CFGINTERRUPTMSIXSENT;
  assign #(out_delay) CFGINTERRUPTMSIXVFENABLE = delay_CFGINTERRUPTMSIXVFENABLE;
  assign #(out_delay) CFGINTERRUPTMSIXVFMASK = delay_CFGINTERRUPTMSIXVFMASK;
  assign #(out_delay) CFGINTERRUPTSENT = delay_CFGINTERRUPTSENT;
  assign #(out_delay) CFGLINKPOWERSTATE = delay_CFGLINKPOWERSTATE;
  assign #(out_delay) CFGLOCALERROR = delay_CFGLOCALERROR;
  assign #(out_delay) CFGLTRENABLE = delay_CFGLTRENABLE;
  assign #(out_delay) CFGLTSSMSTATE = delay_CFGLTSSMSTATE;
  assign #(out_delay) CFGMAXPAYLOAD = delay_CFGMAXPAYLOAD;
  assign #(out_delay) CFGMAXREADREQ = delay_CFGMAXREADREQ;
  assign #(out_delay) CFGMCUPDATEDONE = delay_CFGMCUPDATEDONE;
  assign #(out_delay) CFGMGMTREADDATA = delay_CFGMGMTREADDATA;
  assign #(out_delay) CFGMGMTREADWRITEDONE = delay_CFGMGMTREADWRITEDONE;
  assign #(out_delay) CFGMSGRECEIVED = delay_CFGMSGRECEIVED;
  assign #(out_delay) CFGMSGRECEIVEDDATA = delay_CFGMSGRECEIVEDDATA;
  assign #(out_delay) CFGMSGRECEIVEDTYPE = delay_CFGMSGRECEIVEDTYPE;
  assign #(out_delay) CFGMSGTRANSMITDONE = delay_CFGMSGTRANSMITDONE;
  assign #(out_delay) CFGNEGOTIATEDWIDTH = delay_CFGNEGOTIATEDWIDTH;
  assign #(out_delay) CFGOBFFENABLE = delay_CFGOBFFENABLE;
  assign #(out_delay) CFGPERFUNCSTATUSDATA = delay_CFGPERFUNCSTATUSDATA;
  assign #(out_delay) CFGPERFUNCTIONUPDATEDONE = delay_CFGPERFUNCTIONUPDATEDONE;
  assign #(out_delay) CFGPHYLINKDOWN = delay_CFGPHYLINKDOWN;
  assign #(out_delay) CFGPHYLINKSTATUS = delay_CFGPHYLINKSTATUS;
  assign #(out_delay) CFGPLSTATUSCHANGE = delay_CFGPLSTATUSCHANGE;
  assign #(out_delay) CFGPOWERSTATECHANGEINTERRUPT = delay_CFGPOWERSTATECHANGEINTERRUPT;
  assign #(out_delay) CFGRCBSTATUS = delay_CFGRCBSTATUS;
  assign #(out_delay) CFGTPHFUNCTIONNUM = delay_CFGTPHFUNCTIONNUM;
  assign #(out_delay) CFGTPHREQUESTERENABLE = delay_CFGTPHREQUESTERENABLE;
  assign #(out_delay) CFGTPHSTMODE = delay_CFGTPHSTMODE;
  assign #(out_delay) CFGTPHSTTADDRESS = delay_CFGTPHSTTADDRESS;
  assign #(out_delay) CFGTPHSTTREADENABLE = delay_CFGTPHSTTREADENABLE;
  assign #(out_delay) CFGTPHSTTWRITEBYTEVALID = delay_CFGTPHSTTWRITEBYTEVALID;
  assign #(out_delay) CFGTPHSTTWRITEDATA = delay_CFGTPHSTTWRITEDATA;
  assign #(out_delay) CFGTPHSTTWRITEENABLE = delay_CFGTPHSTTWRITEENABLE;
  assign #(out_delay) CFGVFFLRINPROCESS = delay_CFGVFFLRINPROCESS;
  assign #(out_delay) CFGVFPOWERSTATE = delay_CFGVFPOWERSTATE;
  assign #(out_delay) CFGVFSTATUS = delay_CFGVFSTATUS;
  assign #(out_delay) CFGVFTPHREQUESTERENABLE = delay_CFGVFTPHREQUESTERENABLE;
  assign #(out_delay) CFGVFTPHSTMODE = delay_CFGVFTPHSTMODE;
  assign #(out_delay) DBGDATAOUT = delay_DBGDATAOUT;
  assign #(out_delay) DRPDO = delay_DRPDO;
  assign #(out_delay) DRPRDY = delay_DRPRDY;
  assign #(out_delay) MAXISCQTDATA = delay_MAXISCQTDATA;
  assign #(out_delay) MAXISCQTKEEP = delay_MAXISCQTKEEP;
  assign #(out_delay) MAXISCQTLAST = delay_MAXISCQTLAST;
  assign #(out_delay) MAXISCQTUSER = delay_MAXISCQTUSER;
  assign #(out_delay) MAXISCQTVALID = delay_MAXISCQTVALID;
  assign #(out_delay) MAXISRCTDATA = delay_MAXISRCTDATA;
  assign #(out_delay) MAXISRCTKEEP = delay_MAXISRCTKEEP;
  assign #(out_delay) MAXISRCTLAST = delay_MAXISRCTLAST;
  assign #(out_delay) MAXISRCTUSER = delay_MAXISRCTUSER;
  assign #(out_delay) MAXISRCTVALID = delay_MAXISRCTVALID;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSAL = delay_MICOMPLETIONRAMREADADDRESSAL;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSAU = delay_MICOMPLETIONRAMREADADDRESSAU;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSBL = delay_MICOMPLETIONRAMREADADDRESSBL;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSBU = delay_MICOMPLETIONRAMREADADDRESSBU;
  assign #(out_delay) MICOMPLETIONRAMREADENABLEL = delay_MICOMPLETIONRAMREADENABLEL;
  assign #(out_delay) MICOMPLETIONRAMREADENABLEU = delay_MICOMPLETIONRAMREADENABLEU;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSAL = delay_MICOMPLETIONRAMWRITEADDRESSAL;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSAU = delay_MICOMPLETIONRAMWRITEADDRESSAU;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSBL = delay_MICOMPLETIONRAMWRITEADDRESSBL;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSBU = delay_MICOMPLETIONRAMWRITEADDRESSBU;
  assign #(out_delay) MICOMPLETIONRAMWRITEDATAL = delay_MICOMPLETIONRAMWRITEDATAL;
  assign #(out_delay) MICOMPLETIONRAMWRITEDATAU = delay_MICOMPLETIONRAMWRITEDATAU;
  assign #(out_delay) MICOMPLETIONRAMWRITEENABLEL = delay_MICOMPLETIONRAMWRITEENABLEL;
  assign #(out_delay) MICOMPLETIONRAMWRITEENABLEU = delay_MICOMPLETIONRAMWRITEENABLEU;
  assign #(out_delay) MIREPLAYRAMADDRESS = delay_MIREPLAYRAMADDRESS;
  assign #(out_delay) MIREPLAYRAMREADENABLE = delay_MIREPLAYRAMREADENABLE;
  assign #(out_delay) MIREPLAYRAMWRITEDATA = delay_MIREPLAYRAMWRITEDATA;
  assign #(out_delay) MIREPLAYRAMWRITEENABLE = delay_MIREPLAYRAMWRITEENABLE;
  assign #(out_delay) MIREQUESTRAMREADADDRESSA = delay_MIREQUESTRAMREADADDRESSA;
  assign #(out_delay) MIREQUESTRAMREADADDRESSB = delay_MIREQUESTRAMREADADDRESSB;
  assign #(out_delay) MIREQUESTRAMREADENABLE = delay_MIREQUESTRAMREADENABLE;
  assign #(out_delay) MIREQUESTRAMWRITEADDRESSA = delay_MIREQUESTRAMWRITEADDRESSA;
  assign #(out_delay) MIREQUESTRAMWRITEADDRESSB = delay_MIREQUESTRAMWRITEADDRESSB;
  assign #(out_delay) MIREQUESTRAMWRITEDATA = delay_MIREQUESTRAMWRITEDATA;
  assign #(out_delay) MIREQUESTRAMWRITEENABLE = delay_MIREQUESTRAMWRITEENABLE;
  assign #(out_delay) PCIECQNPREQCOUNT = delay_PCIECQNPREQCOUNT;
  assign #(out_delay) PCIERQSEQNUM = delay_PCIERQSEQNUM;
  assign #(out_delay) PCIERQSEQNUMVLD = delay_PCIERQSEQNUMVLD;
  assign #(out_delay) PCIERQTAG = delay_PCIERQTAG;
  assign #(out_delay) PCIERQTAGAV = delay_PCIERQTAGAV;
  assign #(out_delay) PCIERQTAGVLD = delay_PCIERQTAGVLD;
  assign #(out_delay) PCIETFCNPDAV = delay_PCIETFCNPDAV;
  assign #(out_delay) PCIETFCNPHAV = delay_PCIETFCNPHAV;
  assign #(out_delay) PIPERX0EQCONTROL = delay_PIPERX0EQCONTROL;
  assign #(out_delay) PIPERX0EQLPLFFS = delay_PIPERX0EQLPLFFS;
  assign #(out_delay) PIPERX0EQLPTXPRESET = delay_PIPERX0EQLPTXPRESET;
  assign #(out_delay) PIPERX0EQPRESET = delay_PIPERX0EQPRESET;
  assign #(out_delay) PIPERX0POLARITY = delay_PIPERX0POLARITY;
  assign #(out_delay) PIPERX1EQCONTROL = delay_PIPERX1EQCONTROL;
  assign #(out_delay) PIPERX1EQLPLFFS = delay_PIPERX1EQLPLFFS;
  assign #(out_delay) PIPERX1EQLPTXPRESET = delay_PIPERX1EQLPTXPRESET;
  assign #(out_delay) PIPERX1EQPRESET = delay_PIPERX1EQPRESET;
  assign #(out_delay) PIPERX1POLARITY = delay_PIPERX1POLARITY;
  assign #(out_delay) PIPERX2EQCONTROL = delay_PIPERX2EQCONTROL;
  assign #(out_delay) PIPERX2EQLPLFFS = delay_PIPERX2EQLPLFFS;
  assign #(out_delay) PIPERX2EQLPTXPRESET = delay_PIPERX2EQLPTXPRESET;
  assign #(out_delay) PIPERX2EQPRESET = delay_PIPERX2EQPRESET;
  assign #(out_delay) PIPERX2POLARITY = delay_PIPERX2POLARITY;
  assign #(out_delay) PIPERX3EQCONTROL = delay_PIPERX3EQCONTROL;
  assign #(out_delay) PIPERX3EQLPLFFS = delay_PIPERX3EQLPLFFS;
  assign #(out_delay) PIPERX3EQLPTXPRESET = delay_PIPERX3EQLPTXPRESET;
  assign #(out_delay) PIPERX3EQPRESET = delay_PIPERX3EQPRESET;
  assign #(out_delay) PIPERX3POLARITY = delay_PIPERX3POLARITY;
  assign #(out_delay) PIPERX4EQCONTROL = delay_PIPERX4EQCONTROL;
  assign #(out_delay) PIPERX4EQLPLFFS = delay_PIPERX4EQLPLFFS;
  assign #(out_delay) PIPERX4EQLPTXPRESET = delay_PIPERX4EQLPTXPRESET;
  assign #(out_delay) PIPERX4EQPRESET = delay_PIPERX4EQPRESET;
  assign #(out_delay) PIPERX4POLARITY = delay_PIPERX4POLARITY;
  assign #(out_delay) PIPERX5EQCONTROL = delay_PIPERX5EQCONTROL;
  assign #(out_delay) PIPERX5EQLPLFFS = delay_PIPERX5EQLPLFFS;
  assign #(out_delay) PIPERX5EQLPTXPRESET = delay_PIPERX5EQLPTXPRESET;
  assign #(out_delay) PIPERX5EQPRESET = delay_PIPERX5EQPRESET;
  assign #(out_delay) PIPERX5POLARITY = delay_PIPERX5POLARITY;
  assign #(out_delay) PIPERX6EQCONTROL = delay_PIPERX6EQCONTROL;
  assign #(out_delay) PIPERX6EQLPLFFS = delay_PIPERX6EQLPLFFS;
  assign #(out_delay) PIPERX6EQLPTXPRESET = delay_PIPERX6EQLPTXPRESET;
  assign #(out_delay) PIPERX6EQPRESET = delay_PIPERX6EQPRESET;
  assign #(out_delay) PIPERX6POLARITY = delay_PIPERX6POLARITY;
  assign #(out_delay) PIPERX7EQCONTROL = delay_PIPERX7EQCONTROL;
  assign #(out_delay) PIPERX7EQLPLFFS = delay_PIPERX7EQLPLFFS;
  assign #(out_delay) PIPERX7EQLPTXPRESET = delay_PIPERX7EQLPTXPRESET;
  assign #(out_delay) PIPERX7EQPRESET = delay_PIPERX7EQPRESET;
  assign #(out_delay) PIPERX7POLARITY = delay_PIPERX7POLARITY;
  assign #(out_delay) PIPETX0CHARISK = delay_PIPETX0CHARISK;
  assign #(out_delay) PIPETX0COMPLIANCE = delay_PIPETX0COMPLIANCE;
  assign #(out_delay) PIPETX0DATA = delay_PIPETX0DATA;
  assign #(out_delay) PIPETX0DATAVALID = delay_PIPETX0DATAVALID;
  assign #(out_delay) PIPETX0ELECIDLE = delay_PIPETX0ELECIDLE;
  assign #(out_delay) PIPETX0EQCONTROL = delay_PIPETX0EQCONTROL;
  assign #(out_delay) PIPETX0EQDEEMPH = delay_PIPETX0EQDEEMPH;
  assign #(out_delay) PIPETX0EQPRESET = delay_PIPETX0EQPRESET;
  assign #(out_delay) PIPETX0POWERDOWN = delay_PIPETX0POWERDOWN;
  assign #(out_delay) PIPETX0STARTBLOCK = delay_PIPETX0STARTBLOCK;
  assign #(out_delay) PIPETX0SYNCHEADER = delay_PIPETX0SYNCHEADER;
  assign #(out_delay) PIPETX1CHARISK = delay_PIPETX1CHARISK;
  assign #(out_delay) PIPETX1COMPLIANCE = delay_PIPETX1COMPLIANCE;
  assign #(out_delay) PIPETX1DATA = delay_PIPETX1DATA;
  assign #(out_delay) PIPETX1DATAVALID = delay_PIPETX1DATAVALID;
  assign #(out_delay) PIPETX1ELECIDLE = delay_PIPETX1ELECIDLE;
  assign #(out_delay) PIPETX1EQCONTROL = delay_PIPETX1EQCONTROL;
  assign #(out_delay) PIPETX1EQDEEMPH = delay_PIPETX1EQDEEMPH;
  assign #(out_delay) PIPETX1EQPRESET = delay_PIPETX1EQPRESET;
  assign #(out_delay) PIPETX1POWERDOWN = delay_PIPETX1POWERDOWN;
  assign #(out_delay) PIPETX1STARTBLOCK = delay_PIPETX1STARTBLOCK;
  assign #(out_delay) PIPETX1SYNCHEADER = delay_PIPETX1SYNCHEADER;
  assign #(out_delay) PIPETX2CHARISK = delay_PIPETX2CHARISK;
  assign #(out_delay) PIPETX2COMPLIANCE = delay_PIPETX2COMPLIANCE;
  assign #(out_delay) PIPETX2DATA = delay_PIPETX2DATA;
  assign #(out_delay) PIPETX2DATAVALID = delay_PIPETX2DATAVALID;
  assign #(out_delay) PIPETX2ELECIDLE = delay_PIPETX2ELECIDLE;
  assign #(out_delay) PIPETX2EQCONTROL = delay_PIPETX2EQCONTROL;
  assign #(out_delay) PIPETX2EQDEEMPH = delay_PIPETX2EQDEEMPH;
  assign #(out_delay) PIPETX2EQPRESET = delay_PIPETX2EQPRESET;
  assign #(out_delay) PIPETX2POWERDOWN = delay_PIPETX2POWERDOWN;
  assign #(out_delay) PIPETX2STARTBLOCK = delay_PIPETX2STARTBLOCK;
  assign #(out_delay) PIPETX2SYNCHEADER = delay_PIPETX2SYNCHEADER;
  assign #(out_delay) PIPETX3CHARISK = delay_PIPETX3CHARISK;
  assign #(out_delay) PIPETX3COMPLIANCE = delay_PIPETX3COMPLIANCE;
  assign #(out_delay) PIPETX3DATA = delay_PIPETX3DATA;
  assign #(out_delay) PIPETX3DATAVALID = delay_PIPETX3DATAVALID;
  assign #(out_delay) PIPETX3ELECIDLE = delay_PIPETX3ELECIDLE;
  assign #(out_delay) PIPETX3EQCONTROL = delay_PIPETX3EQCONTROL;
  assign #(out_delay) PIPETX3EQDEEMPH = delay_PIPETX3EQDEEMPH;
  assign #(out_delay) PIPETX3EQPRESET = delay_PIPETX3EQPRESET;
  assign #(out_delay) PIPETX3POWERDOWN = delay_PIPETX3POWERDOWN;
  assign #(out_delay) PIPETX3STARTBLOCK = delay_PIPETX3STARTBLOCK;
  assign #(out_delay) PIPETX3SYNCHEADER = delay_PIPETX3SYNCHEADER;
  assign #(out_delay) PIPETX4CHARISK = delay_PIPETX4CHARISK;
  assign #(out_delay) PIPETX4COMPLIANCE = delay_PIPETX4COMPLIANCE;
  assign #(out_delay) PIPETX4DATA = delay_PIPETX4DATA;
  assign #(out_delay) PIPETX4DATAVALID = delay_PIPETX4DATAVALID;
  assign #(out_delay) PIPETX4ELECIDLE = delay_PIPETX4ELECIDLE;
  assign #(out_delay) PIPETX4EQCONTROL = delay_PIPETX4EQCONTROL;
  assign #(out_delay) PIPETX4EQDEEMPH = delay_PIPETX4EQDEEMPH;
  assign #(out_delay) PIPETX4EQPRESET = delay_PIPETX4EQPRESET;
  assign #(out_delay) PIPETX4POWERDOWN = delay_PIPETX4POWERDOWN;
  assign #(out_delay) PIPETX4STARTBLOCK = delay_PIPETX4STARTBLOCK;
  assign #(out_delay) PIPETX4SYNCHEADER = delay_PIPETX4SYNCHEADER;
  assign #(out_delay) PIPETX5CHARISK = delay_PIPETX5CHARISK;
  assign #(out_delay) PIPETX5COMPLIANCE = delay_PIPETX5COMPLIANCE;
  assign #(out_delay) PIPETX5DATA = delay_PIPETX5DATA;
  assign #(out_delay) PIPETX5DATAVALID = delay_PIPETX5DATAVALID;
  assign #(out_delay) PIPETX5ELECIDLE = delay_PIPETX5ELECIDLE;
  assign #(out_delay) PIPETX5EQCONTROL = delay_PIPETX5EQCONTROL;
  assign #(out_delay) PIPETX5EQDEEMPH = delay_PIPETX5EQDEEMPH;
  assign #(out_delay) PIPETX5EQPRESET = delay_PIPETX5EQPRESET;
  assign #(out_delay) PIPETX5POWERDOWN = delay_PIPETX5POWERDOWN;
  assign #(out_delay) PIPETX5STARTBLOCK = delay_PIPETX5STARTBLOCK;
  assign #(out_delay) PIPETX5SYNCHEADER = delay_PIPETX5SYNCHEADER;
  assign #(out_delay) PIPETX6CHARISK = delay_PIPETX6CHARISK;
  assign #(out_delay) PIPETX6COMPLIANCE = delay_PIPETX6COMPLIANCE;
  assign #(out_delay) PIPETX6DATA = delay_PIPETX6DATA;
  assign #(out_delay) PIPETX6DATAVALID = delay_PIPETX6DATAVALID;
  assign #(out_delay) PIPETX6ELECIDLE = delay_PIPETX6ELECIDLE;
  assign #(out_delay) PIPETX6EQCONTROL = delay_PIPETX6EQCONTROL;
  assign #(out_delay) PIPETX6EQDEEMPH = delay_PIPETX6EQDEEMPH;
  assign #(out_delay) PIPETX6EQPRESET = delay_PIPETX6EQPRESET;
  assign #(out_delay) PIPETX6POWERDOWN = delay_PIPETX6POWERDOWN;
  assign #(out_delay) PIPETX6STARTBLOCK = delay_PIPETX6STARTBLOCK;
  assign #(out_delay) PIPETX6SYNCHEADER = delay_PIPETX6SYNCHEADER;
  assign #(out_delay) PIPETX7CHARISK = delay_PIPETX7CHARISK;
  assign #(out_delay) PIPETX7COMPLIANCE = delay_PIPETX7COMPLIANCE;
  assign #(out_delay) PIPETX7DATA = delay_PIPETX7DATA;
  assign #(out_delay) PIPETX7DATAVALID = delay_PIPETX7DATAVALID;
  assign #(out_delay) PIPETX7ELECIDLE = delay_PIPETX7ELECIDLE;
  assign #(out_delay) PIPETX7EQCONTROL = delay_PIPETX7EQCONTROL;
  assign #(out_delay) PIPETX7EQDEEMPH = delay_PIPETX7EQDEEMPH;
  assign #(out_delay) PIPETX7EQPRESET = delay_PIPETX7EQPRESET;
  assign #(out_delay) PIPETX7POWERDOWN = delay_PIPETX7POWERDOWN;
  assign #(out_delay) PIPETX7STARTBLOCK = delay_PIPETX7STARTBLOCK;
  assign #(out_delay) PIPETX7SYNCHEADER = delay_PIPETX7SYNCHEADER;
  assign #(out_delay) PIPETXDEEMPH = delay_PIPETXDEEMPH;
  assign #(out_delay) PIPETXMARGIN = delay_PIPETXMARGIN;
  assign #(out_delay) PIPETXRATE = delay_PIPETXRATE;
  assign #(out_delay) PIPETXRCVRDET = delay_PIPETXRCVRDET;
  assign #(out_delay) PIPETXRESET = delay_PIPETXRESET;
  assign #(out_delay) PIPETXSWING = delay_PIPETXSWING;
  assign #(out_delay) PLEQINPROGRESS = delay_PLEQINPROGRESS;
  assign #(out_delay) PLEQPHASE = delay_PLEQPHASE;
  assign #(out_delay) PLGEN3PCSRXSLIDE = delay_PLGEN3PCSRXSLIDE;
  assign #(out_delay) SAXISCCTREADY = delay_SAXISCCTREADY;
  assign #(out_delay) SAXISRQTREADY = delay_SAXISRQTREADY;
  
`ifndef XIL_TIMING // unisim
  assign #(INCLK_DELAY) delay_CORECLK = CORECLK;
  assign #(INCLK_DELAY) delay_CORECLKMICOMPLETIONRAML = CORECLKMICOMPLETIONRAML;
  assign #(INCLK_DELAY) delay_CORECLKMICOMPLETIONRAMU = CORECLKMICOMPLETIONRAMU;
  assign #(INCLK_DELAY) delay_CORECLKMIREPLAYRAM = CORECLKMIREPLAYRAM;
  assign #(INCLK_DELAY) delay_CORECLKMIREQUESTRAM = CORECLKMIREQUESTRAM;
  assign #(INCLK_DELAY) delay_DRPCLK = DRPCLK;
  assign #(INCLK_DELAY) delay_PIPECLK = PIPECLK;
  assign #(INCLK_DELAY) delay_RECCLK = RECCLK;
  assign #(INCLK_DELAY) delay_USERCLK = USERCLK;

  assign #(in_delay) delay_CFGCONFIGSPACEENABLE = CFGCONFIGSPACEENABLE;
  assign #(in_delay) delay_CFGDEVID = CFGDEVID;
  assign #(in_delay) delay_CFGDSBUSNUMBER = CFGDSBUSNUMBER;
  assign #(in_delay) delay_CFGDSDEVICENUMBER = CFGDSDEVICENUMBER;
  assign #(in_delay) delay_CFGDSFUNCTIONNUMBER = CFGDSFUNCTIONNUMBER;
  assign #(in_delay) delay_CFGDSN = CFGDSN;
  assign #(in_delay) delay_CFGDSPORTNUMBER = CFGDSPORTNUMBER;
  assign #(in_delay) delay_CFGERRCORIN = CFGERRCORIN;
  assign #(in_delay) delay_CFGERRUNCORIN = CFGERRUNCORIN;
  assign #(in_delay) delay_CFGEXTREADDATA = CFGEXTREADDATA;
  assign #(in_delay) delay_CFGEXTREADDATAVALID = CFGEXTREADDATAVALID;
  assign #(in_delay) delay_CFGFCSEL = CFGFCSEL;
  assign #(in_delay) delay_CFGFLRDONE = CFGFLRDONE;
  assign #(in_delay) delay_CFGHOTRESETIN = CFGHOTRESETIN;
  assign #(in_delay) delay_CFGINPUTUPDATEREQUEST = CFGINPUTUPDATEREQUEST;
  assign #(in_delay) delay_CFGINTERRUPTINT = CFGINTERRUPTINT;
  assign #(in_delay) delay_CFGINTERRUPTMSIATTR = CFGINTERRUPTMSIATTR;
  assign #(in_delay) delay_CFGINTERRUPTMSIFUNCTIONNUMBER = CFGINTERRUPTMSIFUNCTIONNUMBER;
  assign #(in_delay) delay_CFGINTERRUPTMSIINT = CFGINTERRUPTMSIINT;
  assign #(in_delay) delay_CFGINTERRUPTMSIPENDINGSTATUS = CFGINTERRUPTMSIPENDINGSTATUS;
  assign #(in_delay) delay_CFGINTERRUPTMSISELECT = CFGINTERRUPTMSISELECT;
  assign #(in_delay) delay_CFGINTERRUPTMSITPHPRESENT = CFGINTERRUPTMSITPHPRESENT;
  assign #(in_delay) delay_CFGINTERRUPTMSITPHSTTAG = CFGINTERRUPTMSITPHSTTAG;
  assign #(in_delay) delay_CFGINTERRUPTMSITPHTYPE = CFGINTERRUPTMSITPHTYPE;
  assign #(in_delay) delay_CFGINTERRUPTMSIXADDRESS = CFGINTERRUPTMSIXADDRESS;
  assign #(in_delay) delay_CFGINTERRUPTMSIXDATA = CFGINTERRUPTMSIXDATA;
  assign #(in_delay) delay_CFGINTERRUPTMSIXINT = CFGINTERRUPTMSIXINT;
  assign #(in_delay) delay_CFGINTERRUPTPENDING = CFGINTERRUPTPENDING;
  assign #(in_delay) delay_CFGLINKTRAININGENABLE = CFGLINKTRAININGENABLE;
  assign #(in_delay) delay_CFGMCUPDATEREQUEST = CFGMCUPDATEREQUEST;
  assign #(in_delay) delay_CFGMGMTADDR = CFGMGMTADDR;
  assign #(in_delay) delay_CFGMGMTBYTEENABLE = CFGMGMTBYTEENABLE;
  assign #(in_delay) delay_CFGMGMTREAD = CFGMGMTREAD;
  assign #(in_delay) delay_CFGMGMTTYPE1CFGREGACCESS = CFGMGMTTYPE1CFGREGACCESS;
  assign #(in_delay) delay_CFGMGMTWRITE = CFGMGMTWRITE;
  assign #(in_delay) delay_CFGMGMTWRITEDATA = CFGMGMTWRITEDATA;
  assign #(in_delay) delay_CFGMSGTRANSMIT = CFGMSGTRANSMIT;
  assign #(in_delay) delay_CFGMSGTRANSMITDATA = CFGMSGTRANSMITDATA;
  assign #(in_delay) delay_CFGMSGTRANSMITTYPE = CFGMSGTRANSMITTYPE;
  assign #(in_delay) delay_CFGPERFUNCSTATUSCONTROL = CFGPERFUNCSTATUSCONTROL;
  assign #(in_delay) delay_CFGPERFUNCTIONNUMBER = CFGPERFUNCTIONNUMBER;
  assign #(in_delay) delay_CFGPERFUNCTIONOUTPUTREQUEST = CFGPERFUNCTIONOUTPUTREQUEST;
  assign #(in_delay) delay_CFGPOWERSTATECHANGEACK = CFGPOWERSTATECHANGEACK;
  assign #(in_delay) delay_CFGREQPMTRANSITIONL23READY = CFGREQPMTRANSITIONL23READY;
  assign #(in_delay) delay_CFGREVID = CFGREVID;
  assign #(in_delay) delay_CFGSUBSYSID = CFGSUBSYSID;
  assign #(in_delay) delay_CFGSUBSYSVENDID = CFGSUBSYSVENDID;
  assign #(in_delay) delay_CFGTPHSTTREADDATA = CFGTPHSTTREADDATA;
  assign #(in_delay) delay_CFGTPHSTTREADDATAVALID = CFGTPHSTTREADDATAVALID;
  assign #(in_delay) delay_CFGVENDID = CFGVENDID;
  assign #(in_delay) delay_CFGVFFLRDONE = CFGVFFLRDONE;
  assign #(in_delay) delay_DRPADDR = DRPADDR;
  assign #(in_delay) delay_DRPDI = DRPDI;
  assign #(in_delay) delay_DRPEN = DRPEN;
  assign #(in_delay) delay_DRPWE = DRPWE;
  assign #(in_delay) delay_MAXISCQTREADY = MAXISCQTREADY;
  assign #(in_delay) delay_MAXISRCTREADY = MAXISRCTREADY;
  assign #(in_delay) delay_MGMTRESETN = MGMTRESETN;
  assign #(in_delay) delay_MGMTSTICKYRESETN = MGMTSTICKYRESETN;
  assign #(in_delay) delay_MICOMPLETIONRAMREADDATA = MICOMPLETIONRAMREADDATA;
  assign #(in_delay) delay_MIREPLAYRAMREADDATA = MIREPLAYRAMREADDATA;
  assign #(in_delay) delay_MIREQUESTRAMREADDATA = MIREQUESTRAMREADDATA;
  assign #(in_delay) delay_PCIECQNPREQ = PCIECQNPREQ;
  assign #(in_delay) delay_PIPEEQFS = PIPEEQFS;
  assign #(in_delay) delay_PIPEEQLF = PIPEEQLF;
  assign #(in_delay) delay_PIPERESETN = PIPERESETN;
  assign #(in_delay) delay_PIPERX0CHARISK = PIPERX0CHARISK;
  assign #(in_delay) delay_PIPERX0DATA = PIPERX0DATA;
  assign #(in_delay) delay_PIPERX0DATAVALID = PIPERX0DATAVALID;
  assign #(in_delay) delay_PIPERX0ELECIDLE = PIPERX0ELECIDLE;
  assign #(in_delay) delay_PIPERX0EQDONE = PIPERX0EQDONE;
  assign #(in_delay) delay_PIPERX0EQLPADAPTDONE = PIPERX0EQLPADAPTDONE;
  assign #(in_delay) delay_PIPERX0EQLPLFFSSEL = PIPERX0EQLPLFFSSEL;
  assign #(in_delay) delay_PIPERX0EQLPNEWTXCOEFFORPRESET = PIPERX0EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) delay_PIPERX0PHYSTATUS = PIPERX0PHYSTATUS;
  assign #(in_delay) delay_PIPERX0STARTBLOCK = PIPERX0STARTBLOCK;
  assign #(in_delay) delay_PIPERX0STATUS = PIPERX0STATUS;
  assign #(in_delay) delay_PIPERX0SYNCHEADER = PIPERX0SYNCHEADER;
  assign #(in_delay) delay_PIPERX0VALID = PIPERX0VALID;
  assign #(in_delay) delay_PIPERX1CHARISK = PIPERX1CHARISK;
  assign #(in_delay) delay_PIPERX1DATA = PIPERX1DATA;
  assign #(in_delay) delay_PIPERX1DATAVALID = PIPERX1DATAVALID;
  assign #(in_delay) delay_PIPERX1ELECIDLE = PIPERX1ELECIDLE;
  assign #(in_delay) delay_PIPERX1EQDONE = PIPERX1EQDONE;
  assign #(in_delay) delay_PIPERX1EQLPADAPTDONE = PIPERX1EQLPADAPTDONE;
  assign #(in_delay) delay_PIPERX1EQLPLFFSSEL = PIPERX1EQLPLFFSSEL;
  assign #(in_delay) delay_PIPERX1EQLPNEWTXCOEFFORPRESET = PIPERX1EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) delay_PIPERX1PHYSTATUS = PIPERX1PHYSTATUS;
  assign #(in_delay) delay_PIPERX1STARTBLOCK = PIPERX1STARTBLOCK;
  assign #(in_delay) delay_PIPERX1STATUS = PIPERX1STATUS;
  assign #(in_delay) delay_PIPERX1SYNCHEADER = PIPERX1SYNCHEADER;
  assign #(in_delay) delay_PIPERX1VALID = PIPERX1VALID;
  assign #(in_delay) delay_PIPERX2CHARISK = PIPERX2CHARISK;
  assign #(in_delay) delay_PIPERX2DATA = PIPERX2DATA;
  assign #(in_delay) delay_PIPERX2DATAVALID = PIPERX2DATAVALID;
  assign #(in_delay) delay_PIPERX2ELECIDLE = PIPERX2ELECIDLE;
  assign #(in_delay) delay_PIPERX2EQDONE = PIPERX2EQDONE;
  assign #(in_delay) delay_PIPERX2EQLPADAPTDONE = PIPERX2EQLPADAPTDONE;
  assign #(in_delay) delay_PIPERX2EQLPLFFSSEL = PIPERX2EQLPLFFSSEL;
  assign #(in_delay) delay_PIPERX2EQLPNEWTXCOEFFORPRESET = PIPERX2EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) delay_PIPERX2PHYSTATUS = PIPERX2PHYSTATUS;
  assign #(in_delay) delay_PIPERX2STARTBLOCK = PIPERX2STARTBLOCK;
  assign #(in_delay) delay_PIPERX2STATUS = PIPERX2STATUS;
  assign #(in_delay) delay_PIPERX2SYNCHEADER = PIPERX2SYNCHEADER;
  assign #(in_delay) delay_PIPERX2VALID = PIPERX2VALID;
  assign #(in_delay) delay_PIPERX3CHARISK = PIPERX3CHARISK;
  assign #(in_delay) delay_PIPERX3DATA = PIPERX3DATA;
  assign #(in_delay) delay_PIPERX3DATAVALID = PIPERX3DATAVALID;
  assign #(in_delay) delay_PIPERX3ELECIDLE = PIPERX3ELECIDLE;
  assign #(in_delay) delay_PIPERX3EQDONE = PIPERX3EQDONE;
  assign #(in_delay) delay_PIPERX3EQLPADAPTDONE = PIPERX3EQLPADAPTDONE;
  assign #(in_delay) delay_PIPERX3EQLPLFFSSEL = PIPERX3EQLPLFFSSEL;
  assign #(in_delay) delay_PIPERX3EQLPNEWTXCOEFFORPRESET = PIPERX3EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) delay_PIPERX3PHYSTATUS = PIPERX3PHYSTATUS;
  assign #(in_delay) delay_PIPERX3STARTBLOCK = PIPERX3STARTBLOCK;
  assign #(in_delay) delay_PIPERX3STATUS = PIPERX3STATUS;
  assign #(in_delay) delay_PIPERX3SYNCHEADER = PIPERX3SYNCHEADER;
  assign #(in_delay) delay_PIPERX3VALID = PIPERX3VALID;
  assign #(in_delay) delay_PIPERX4CHARISK = PIPERX4CHARISK;
  assign #(in_delay) delay_PIPERX4DATA = PIPERX4DATA;
  assign #(in_delay) delay_PIPERX4DATAVALID = PIPERX4DATAVALID;
  assign #(in_delay) delay_PIPERX4ELECIDLE = PIPERX4ELECIDLE;
  assign #(in_delay) delay_PIPERX4EQDONE = PIPERX4EQDONE;
  assign #(in_delay) delay_PIPERX4EQLPADAPTDONE = PIPERX4EQLPADAPTDONE;
  assign #(in_delay) delay_PIPERX4EQLPLFFSSEL = PIPERX4EQLPLFFSSEL;
  assign #(in_delay) delay_PIPERX4EQLPNEWTXCOEFFORPRESET = PIPERX4EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) delay_PIPERX4PHYSTATUS = PIPERX4PHYSTATUS;
  assign #(in_delay) delay_PIPERX4STARTBLOCK = PIPERX4STARTBLOCK;
  assign #(in_delay) delay_PIPERX4STATUS = PIPERX4STATUS;
  assign #(in_delay) delay_PIPERX4SYNCHEADER = PIPERX4SYNCHEADER;
  assign #(in_delay) delay_PIPERX4VALID = PIPERX4VALID;
  assign #(in_delay) delay_PIPERX5CHARISK = PIPERX5CHARISK;
  assign #(in_delay) delay_PIPERX5DATA = PIPERX5DATA;
  assign #(in_delay) delay_PIPERX5DATAVALID = PIPERX5DATAVALID;
  assign #(in_delay) delay_PIPERX5ELECIDLE = PIPERX5ELECIDLE;
  assign #(in_delay) delay_PIPERX5EQDONE = PIPERX5EQDONE;
  assign #(in_delay) delay_PIPERX5EQLPADAPTDONE = PIPERX5EQLPADAPTDONE;
  assign #(in_delay) delay_PIPERX5EQLPLFFSSEL = PIPERX5EQLPLFFSSEL;
  assign #(in_delay) delay_PIPERX5EQLPNEWTXCOEFFORPRESET = PIPERX5EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) delay_PIPERX5PHYSTATUS = PIPERX5PHYSTATUS;
  assign #(in_delay) delay_PIPERX5STARTBLOCK = PIPERX5STARTBLOCK;
  assign #(in_delay) delay_PIPERX5STATUS = PIPERX5STATUS;
  assign #(in_delay) delay_PIPERX5SYNCHEADER = PIPERX5SYNCHEADER;
  assign #(in_delay) delay_PIPERX5VALID = PIPERX5VALID;
  assign #(in_delay) delay_PIPERX6CHARISK = PIPERX6CHARISK;
  assign #(in_delay) delay_PIPERX6DATA = PIPERX6DATA;
  assign #(in_delay) delay_PIPERX6DATAVALID = PIPERX6DATAVALID;
  assign #(in_delay) delay_PIPERX6ELECIDLE = PIPERX6ELECIDLE;
  assign #(in_delay) delay_PIPERX6EQDONE = PIPERX6EQDONE;
  assign #(in_delay) delay_PIPERX6EQLPADAPTDONE = PIPERX6EQLPADAPTDONE;
  assign #(in_delay) delay_PIPERX6EQLPLFFSSEL = PIPERX6EQLPLFFSSEL;
  assign #(in_delay) delay_PIPERX6EQLPNEWTXCOEFFORPRESET = PIPERX6EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) delay_PIPERX6PHYSTATUS = PIPERX6PHYSTATUS;
  assign #(in_delay) delay_PIPERX6STARTBLOCK = PIPERX6STARTBLOCK;
  assign #(in_delay) delay_PIPERX6STATUS = PIPERX6STATUS;
  assign #(in_delay) delay_PIPERX6SYNCHEADER = PIPERX6SYNCHEADER;
  assign #(in_delay) delay_PIPERX6VALID = PIPERX6VALID;
  assign #(in_delay) delay_PIPERX7CHARISK = PIPERX7CHARISK;
  assign #(in_delay) delay_PIPERX7DATA = PIPERX7DATA;
  assign #(in_delay) delay_PIPERX7DATAVALID = PIPERX7DATAVALID;
  assign #(in_delay) delay_PIPERX7ELECIDLE = PIPERX7ELECIDLE;
  assign #(in_delay) delay_PIPERX7EQDONE = PIPERX7EQDONE;
  assign #(in_delay) delay_PIPERX7EQLPADAPTDONE = PIPERX7EQLPADAPTDONE;
  assign #(in_delay) delay_PIPERX7EQLPLFFSSEL = PIPERX7EQLPLFFSSEL;
  assign #(in_delay) delay_PIPERX7EQLPNEWTXCOEFFORPRESET = PIPERX7EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) delay_PIPERX7PHYSTATUS = PIPERX7PHYSTATUS;
  assign #(in_delay) delay_PIPERX7STARTBLOCK = PIPERX7STARTBLOCK;
  assign #(in_delay) delay_PIPERX7STATUS = PIPERX7STATUS;
  assign #(in_delay) delay_PIPERX7SYNCHEADER = PIPERX7SYNCHEADER;
  assign #(in_delay) delay_PIPERX7VALID = PIPERX7VALID;
  assign #(in_delay) delay_PIPETX0EQCOEFF = PIPETX0EQCOEFF;
  assign #(in_delay) delay_PIPETX0EQDONE = PIPETX0EQDONE;
  assign #(in_delay) delay_PIPETX1EQCOEFF = PIPETX1EQCOEFF;
  assign #(in_delay) delay_PIPETX1EQDONE = PIPETX1EQDONE;
  assign #(in_delay) delay_PIPETX2EQCOEFF = PIPETX2EQCOEFF;
  assign #(in_delay) delay_PIPETX2EQDONE = PIPETX2EQDONE;
  assign #(in_delay) delay_PIPETX3EQCOEFF = PIPETX3EQCOEFF;
  assign #(in_delay) delay_PIPETX3EQDONE = PIPETX3EQDONE;
  assign #(in_delay) delay_PIPETX4EQCOEFF = PIPETX4EQCOEFF;
  assign #(in_delay) delay_PIPETX4EQDONE = PIPETX4EQDONE;
  assign #(in_delay) delay_PIPETX5EQCOEFF = PIPETX5EQCOEFF;
  assign #(in_delay) delay_PIPETX5EQDONE = PIPETX5EQDONE;
  assign #(in_delay) delay_PIPETX6EQCOEFF = PIPETX6EQCOEFF;
  assign #(in_delay) delay_PIPETX6EQDONE = PIPETX6EQDONE;
  assign #(in_delay) delay_PIPETX7EQCOEFF = PIPETX7EQCOEFF;
  assign #(in_delay) delay_PIPETX7EQDONE = PIPETX7EQDONE;
  assign #(in_delay) delay_PLDISABLESCRAMBLER = PLDISABLESCRAMBLER;
  assign #(in_delay) delay_PLEQRESETEIEOSCOUNT = PLEQRESETEIEOSCOUNT;
  assign #(in_delay) delay_PLGEN3PCSDISABLE = PLGEN3PCSDISABLE;
  assign #(in_delay) delay_PLGEN3PCSRXSYNCDONE = PLGEN3PCSRXSYNCDONE;
  assign #(in_delay) delay_RESETN = RESETN;
  assign #(in_delay) delay_SAXISCCTDATA = SAXISCCTDATA;
  assign #(in_delay) delay_SAXISCCTKEEP = SAXISCCTKEEP;
  assign #(in_delay) delay_SAXISCCTLAST = SAXISCCTLAST;
  assign #(in_delay) delay_SAXISCCTUSER = SAXISCCTUSER;
  assign #(in_delay) delay_SAXISCCTVALID = SAXISCCTVALID;
  assign #(in_delay) delay_SAXISRQTDATA = SAXISRQTDATA;
  assign #(in_delay) delay_SAXISRQTKEEP = SAXISRQTKEEP;
  assign #(in_delay) delay_SAXISRQTLAST = SAXISRQTLAST;
  assign #(in_delay) delay_SAXISRQTUSER = SAXISRQTUSER;
  assign #(in_delay) delay_SAXISRQTVALID = SAXISRQTVALID;
`endif //  `ifndef XIL_TIMING

`ifdef XIL_TIMING //Simprim
  assign delay_CORECLKMICOMPLETIONRAML = CORECLKMICOMPLETIONRAML;
  assign delay_CORECLKMICOMPLETIONRAMU = CORECLKMICOMPLETIONRAMU;
  assign delay_CORECLKMIREPLAYRAM = CORECLKMIREPLAYRAM;
  assign delay_CORECLKMIREQUESTRAM = CORECLKMIREQUESTRAM;
  assign delay_MGMTRESETN = MGMTRESETN;
  assign delay_MGMTSTICKYRESETN = MGMTSTICKYRESETN;
  assign delay_PIPERESETN = PIPERESETN;
  assign delay_RESETN = RESETN;
`endif

  B_PCIE_3_0 #(
    .ARI_CAP_ENABLE (ARI_CAP_ENABLE),
    .AXISTEN_IF_CC_ALIGNMENT_MODE (AXISTEN_IF_CC_ALIGNMENT_MODE),
    .AXISTEN_IF_CC_PARITY_CHK (AXISTEN_IF_CC_PARITY_CHK),
    .AXISTEN_IF_CQ_ALIGNMENT_MODE (AXISTEN_IF_CQ_ALIGNMENT_MODE),
    .AXISTEN_IF_ENABLE_CLIENT_TAG (AXISTEN_IF_ENABLE_CLIENT_TAG),
    .AXISTEN_IF_ENABLE_MSG_ROUTE (AXISTEN_IF_ENABLE_MSG_ROUTE),
    .AXISTEN_IF_ENABLE_RX_MSG_INTFC (AXISTEN_IF_ENABLE_RX_MSG_INTFC),
    .AXISTEN_IF_RC_ALIGNMENT_MODE (AXISTEN_IF_RC_ALIGNMENT_MODE),
    .AXISTEN_IF_RC_STRADDLE (AXISTEN_IF_RC_STRADDLE),
    .AXISTEN_IF_RQ_ALIGNMENT_MODE (AXISTEN_IF_RQ_ALIGNMENT_MODE),
    .AXISTEN_IF_RQ_PARITY_CHK (AXISTEN_IF_RQ_PARITY_CHK),
    .AXISTEN_IF_WIDTH (AXISTEN_IF_WIDTH),
    .CRM_CORE_CLK_FREQ_500 (CRM_CORE_CLK_FREQ_500),
    .CRM_USER_CLK_FREQ (CRM_USER_CLK_FREQ),
    .DNSTREAM_LINK_NUM (DNSTREAM_LINK_NUM),
    .GEN3_PCS_AUTO_REALIGN (GEN3_PCS_AUTO_REALIGN),
    .GEN3_PCS_RX_ELECIDLE_INTERNAL (GEN3_PCS_RX_ELECIDLE_INTERNAL),
    .LL_ACK_TIMEOUT (LL_ACK_TIMEOUT),
    .LL_ACK_TIMEOUT_EN (LL_ACK_TIMEOUT_EN),
    .LL_ACK_TIMEOUT_FUNC (LL_ACK_TIMEOUT_FUNC),
    .LL_CPL_FC_UPDATE_TIMER (LL_CPL_FC_UPDATE_TIMER),
    .LL_CPL_FC_UPDATE_TIMER_OVERRIDE (LL_CPL_FC_UPDATE_TIMER_OVERRIDE),
    .LL_FC_UPDATE_TIMER (LL_FC_UPDATE_TIMER),
    .LL_FC_UPDATE_TIMER_OVERRIDE (LL_FC_UPDATE_TIMER_OVERRIDE),
    .LL_NP_FC_UPDATE_TIMER (LL_NP_FC_UPDATE_TIMER),
    .LL_NP_FC_UPDATE_TIMER_OVERRIDE (LL_NP_FC_UPDATE_TIMER_OVERRIDE),
    .LL_P_FC_UPDATE_TIMER (LL_P_FC_UPDATE_TIMER),
    .LL_P_FC_UPDATE_TIMER_OVERRIDE (LL_P_FC_UPDATE_TIMER_OVERRIDE),
    .LL_REPLAY_TIMEOUT (LL_REPLAY_TIMEOUT),
    .LL_REPLAY_TIMEOUT_EN (LL_REPLAY_TIMEOUT_EN),
    .LL_REPLAY_TIMEOUT_FUNC (LL_REPLAY_TIMEOUT_FUNC),
    .LTR_TX_MESSAGE_MINIMUM_INTERVAL (LTR_TX_MESSAGE_MINIMUM_INTERVAL),
    .LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE (LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE),
    .LTR_TX_MESSAGE_ON_LTR_ENABLE (LTR_TX_MESSAGE_ON_LTR_ENABLE),
    .PF0_AER_CAP_ECRC_CHECK_CAPABLE (PF0_AER_CAP_ECRC_CHECK_CAPABLE),
    .PF0_AER_CAP_ECRC_GEN_CAPABLE (PF0_AER_CAP_ECRC_GEN_CAPABLE),
    .PF0_AER_CAP_NEXTPTR (PF0_AER_CAP_NEXTPTR),
    .PF0_ARI_CAP_NEXTPTR (PF0_ARI_CAP_NEXTPTR),
    .PF0_ARI_CAP_NEXT_FUNC (PF0_ARI_CAP_NEXT_FUNC),
    .PF0_ARI_CAP_VER (PF0_ARI_CAP_VER),
    .PF0_BAR0_APERTURE_SIZE (PF0_BAR0_APERTURE_SIZE),
    .PF0_BAR0_CONTROL (PF0_BAR0_CONTROL),
    .PF0_BAR1_APERTURE_SIZE (PF0_BAR1_APERTURE_SIZE),
    .PF0_BAR1_CONTROL (PF0_BAR1_CONTROL),
    .PF0_BAR2_APERTURE_SIZE (PF0_BAR2_APERTURE_SIZE),
    .PF0_BAR2_CONTROL (PF0_BAR2_CONTROL),
    .PF0_BAR3_APERTURE_SIZE (PF0_BAR3_APERTURE_SIZE),
    .PF0_BAR3_CONTROL (PF0_BAR3_CONTROL),
    .PF0_BAR4_APERTURE_SIZE (PF0_BAR4_APERTURE_SIZE),
    .PF0_BAR4_CONTROL (PF0_BAR4_CONTROL),
    .PF0_BAR5_APERTURE_SIZE (PF0_BAR5_APERTURE_SIZE),
    .PF0_BAR5_CONTROL (PF0_BAR5_CONTROL),
    .PF0_BIST_REGISTER (PF0_BIST_REGISTER),
    .PF0_CAPABILITY_POINTER (PF0_CAPABILITY_POINTER),
    .PF0_CLASS_CODE (PF0_CLASS_CODE),
    .PF0_DEVICE_ID (PF0_DEVICE_ID),
    .PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT (PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT),
    .PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT (PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT),
    .PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT (PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT),
    .PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE (PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE),
    .PF0_DEV_CAP2_LTR_SUPPORT (PF0_DEV_CAP2_LTR_SUPPORT),
    .PF0_DEV_CAP2_OBFF_SUPPORT (PF0_DEV_CAP2_OBFF_SUPPORT),
    .PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT (PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT),
    .PF0_DEV_CAP_ENDPOINT_L0S_LATENCY (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY),
    .PF0_DEV_CAP_ENDPOINT_L1_LATENCY (PF0_DEV_CAP_ENDPOINT_L1_LATENCY),
    .PF0_DEV_CAP_EXT_TAG_SUPPORTED (PF0_DEV_CAP_EXT_TAG_SUPPORTED),
    .PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE (PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE),
    .PF0_DEV_CAP_MAX_PAYLOAD_SIZE (PF0_DEV_CAP_MAX_PAYLOAD_SIZE),
    .PF0_DPA_CAP_NEXTPTR (PF0_DPA_CAP_NEXTPTR),
    .PF0_DPA_CAP_SUB_STATE_CONTROL (PF0_DPA_CAP_SUB_STATE_CONTROL),
    .PF0_DPA_CAP_SUB_STATE_CONTROL_EN (PF0_DPA_CAP_SUB_STATE_CONTROL_EN),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7),
    .PF0_DPA_CAP_VER (PF0_DPA_CAP_VER),
    .PF0_DSN_CAP_NEXTPTR (PF0_DSN_CAP_NEXTPTR),
    .PF0_EXPANSION_ROM_APERTURE_SIZE (PF0_EXPANSION_ROM_APERTURE_SIZE),
    .PF0_EXPANSION_ROM_ENABLE (PF0_EXPANSION_ROM_ENABLE),
    .PF0_INTERRUPT_LINE (PF0_INTERRUPT_LINE),
    .PF0_INTERRUPT_PIN (PF0_INTERRUPT_PIN),
    .PF0_LINK_CAP_ASPM_SUPPORT (PF0_LINK_CAP_ASPM_SUPPORT),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3),
    .PF0_LINK_STATUS_SLOT_CLOCK_CONFIG (PF0_LINK_STATUS_SLOT_CLOCK_CONFIG),
    .PF0_LTR_CAP_MAX_NOSNOOP_LAT (PF0_LTR_CAP_MAX_NOSNOOP_LAT),
    .PF0_LTR_CAP_MAX_SNOOP_LAT (PF0_LTR_CAP_MAX_SNOOP_LAT),
    .PF0_LTR_CAP_NEXTPTR (PF0_LTR_CAP_NEXTPTR),
    .PF0_LTR_CAP_VER (PF0_LTR_CAP_VER),
    .PF0_MSIX_CAP_NEXTPTR (PF0_MSIX_CAP_NEXTPTR),
    .PF0_MSIX_CAP_PBA_BIR (PF0_MSIX_CAP_PBA_BIR),
    .PF0_MSIX_CAP_PBA_OFFSET (PF0_MSIX_CAP_PBA_OFFSET),
    .PF0_MSIX_CAP_TABLE_BIR (PF0_MSIX_CAP_TABLE_BIR),
    .PF0_MSIX_CAP_TABLE_OFFSET (PF0_MSIX_CAP_TABLE_OFFSET),
    .PF0_MSIX_CAP_TABLE_SIZE (PF0_MSIX_CAP_TABLE_SIZE),
    .PF0_MSI_CAP_MULTIMSGCAP (PF0_MSI_CAP_MULTIMSGCAP),
    .PF0_MSI_CAP_NEXTPTR (PF0_MSI_CAP_NEXTPTR),
    .PF0_PB_CAP_NEXTPTR (PF0_PB_CAP_NEXTPTR),
    .PF0_PB_CAP_SYSTEM_ALLOCATED (PF0_PB_CAP_SYSTEM_ALLOCATED),
    .PF0_PB_CAP_VER (PF0_PB_CAP_VER),
    .PF0_PM_CAP_ID (PF0_PM_CAP_ID),
    .PF0_PM_CAP_NEXTPTR (PF0_PM_CAP_NEXTPTR),
    .PF0_PM_CAP_PMESUPPORT_D0 (PF0_PM_CAP_PMESUPPORT_D0),
    .PF0_PM_CAP_PMESUPPORT_D1 (PF0_PM_CAP_PMESUPPORT_D1),
    .PF0_PM_CAP_PMESUPPORT_D3HOT (PF0_PM_CAP_PMESUPPORT_D3HOT),
    .PF0_PM_CAP_SUPP_D1_STATE (PF0_PM_CAP_SUPP_D1_STATE),
    .PF0_PM_CAP_VER_ID (PF0_PM_CAP_VER_ID),
    .PF0_PM_CSR_NOSOFTRESET (PF0_PM_CSR_NOSOFTRESET),
    .PF0_RBAR_CAP_ENABLE (PF0_RBAR_CAP_ENABLE),
    .PF0_RBAR_CAP_INDEX0 (PF0_RBAR_CAP_INDEX0),
    .PF0_RBAR_CAP_INDEX1 (PF0_RBAR_CAP_INDEX1),
    .PF0_RBAR_CAP_INDEX2 (PF0_RBAR_CAP_INDEX2),
    .PF0_RBAR_CAP_NEXTPTR (PF0_RBAR_CAP_NEXTPTR),
    .PF0_RBAR_CAP_SIZE0 (PF0_RBAR_CAP_SIZE0),
    .PF0_RBAR_CAP_SIZE1 (PF0_RBAR_CAP_SIZE1),
    .PF0_RBAR_CAP_SIZE2 (PF0_RBAR_CAP_SIZE2),
    .PF0_RBAR_CAP_VER (PF0_RBAR_CAP_VER),
    .PF0_RBAR_NUM (PF0_RBAR_NUM),
    .PF0_REVISION_ID (PF0_REVISION_ID),
    .PF0_SRIOV_BAR0_APERTURE_SIZE (PF0_SRIOV_BAR0_APERTURE_SIZE),
    .PF0_SRIOV_BAR0_CONTROL (PF0_SRIOV_BAR0_CONTROL),
    .PF0_SRIOV_BAR1_APERTURE_SIZE (PF0_SRIOV_BAR1_APERTURE_SIZE),
    .PF0_SRIOV_BAR1_CONTROL (PF0_SRIOV_BAR1_CONTROL),
    .PF0_SRIOV_BAR2_APERTURE_SIZE (PF0_SRIOV_BAR2_APERTURE_SIZE),
    .PF0_SRIOV_BAR2_CONTROL (PF0_SRIOV_BAR2_CONTROL),
    .PF0_SRIOV_BAR3_APERTURE_SIZE (PF0_SRIOV_BAR3_APERTURE_SIZE),
    .PF0_SRIOV_BAR3_CONTROL (PF0_SRIOV_BAR3_CONTROL),
    .PF0_SRIOV_BAR4_APERTURE_SIZE (PF0_SRIOV_BAR4_APERTURE_SIZE),
    .PF0_SRIOV_BAR4_CONTROL (PF0_SRIOV_BAR4_CONTROL),
    .PF0_SRIOV_BAR5_APERTURE_SIZE (PF0_SRIOV_BAR5_APERTURE_SIZE),
    .PF0_SRIOV_BAR5_CONTROL (PF0_SRIOV_BAR5_CONTROL),
    .PF0_SRIOV_CAP_INITIAL_VF (PF0_SRIOV_CAP_INITIAL_VF),
    .PF0_SRIOV_CAP_NEXTPTR (PF0_SRIOV_CAP_NEXTPTR),
    .PF0_SRIOV_CAP_TOTAL_VF (PF0_SRIOV_CAP_TOTAL_VF),
    .PF0_SRIOV_CAP_VER (PF0_SRIOV_CAP_VER),
    .PF0_SRIOV_FIRST_VF_OFFSET (PF0_SRIOV_FIRST_VF_OFFSET),
    .PF0_SRIOV_FUNC_DEP_LINK (PF0_SRIOV_FUNC_DEP_LINK),
    .PF0_SRIOV_SUPPORTED_PAGE_SIZE (PF0_SRIOV_SUPPORTED_PAGE_SIZE),
    .PF0_SRIOV_VF_DEVICE_ID (PF0_SRIOV_VF_DEVICE_ID),
    .PF0_SUBSYSTEM_ID (PF0_SUBSYSTEM_ID),
    .PF0_TPHR_CAP_DEV_SPECIFIC_MODE (PF0_TPHR_CAP_DEV_SPECIFIC_MODE),
    .PF0_TPHR_CAP_ENABLE (PF0_TPHR_CAP_ENABLE),
    .PF0_TPHR_CAP_INT_VEC_MODE (PF0_TPHR_CAP_INT_VEC_MODE),
    .PF0_TPHR_CAP_NEXTPTR (PF0_TPHR_CAP_NEXTPTR),
    .PF0_TPHR_CAP_ST_MODE_SEL (PF0_TPHR_CAP_ST_MODE_SEL),
    .PF0_TPHR_CAP_ST_TABLE_LOC (PF0_TPHR_CAP_ST_TABLE_LOC),
    .PF0_TPHR_CAP_ST_TABLE_SIZE (PF0_TPHR_CAP_ST_TABLE_SIZE),
    .PF0_TPHR_CAP_VER (PF0_TPHR_CAP_VER),
    .PF0_VC_CAP_NEXTPTR (PF0_VC_CAP_NEXTPTR),
    .PF0_VC_CAP_VER (PF0_VC_CAP_VER),
    .PF1_AER_CAP_ECRC_CHECK_CAPABLE (PF1_AER_CAP_ECRC_CHECK_CAPABLE),
    .PF1_AER_CAP_ECRC_GEN_CAPABLE (PF1_AER_CAP_ECRC_GEN_CAPABLE),
    .PF1_AER_CAP_NEXTPTR (PF1_AER_CAP_NEXTPTR),
    .PF1_ARI_CAP_NEXTPTR (PF1_ARI_CAP_NEXTPTR),
    .PF1_ARI_CAP_NEXT_FUNC (PF1_ARI_CAP_NEXT_FUNC),
    .PF1_BAR0_APERTURE_SIZE (PF1_BAR0_APERTURE_SIZE),
    .PF1_BAR0_CONTROL (PF1_BAR0_CONTROL),
    .PF1_BAR1_APERTURE_SIZE (PF1_BAR1_APERTURE_SIZE),
    .PF1_BAR1_CONTROL (PF1_BAR1_CONTROL),
    .PF1_BAR2_APERTURE_SIZE (PF1_BAR2_APERTURE_SIZE),
    .PF1_BAR2_CONTROL (PF1_BAR2_CONTROL),
    .PF1_BAR3_APERTURE_SIZE (PF1_BAR3_APERTURE_SIZE),
    .PF1_BAR3_CONTROL (PF1_BAR3_CONTROL),
    .PF1_BAR4_APERTURE_SIZE (PF1_BAR4_APERTURE_SIZE),
    .PF1_BAR4_CONTROL (PF1_BAR4_CONTROL),
    .PF1_BAR5_APERTURE_SIZE (PF1_BAR5_APERTURE_SIZE),
    .PF1_BAR5_CONTROL (PF1_BAR5_CONTROL),
    .PF1_BIST_REGISTER (PF1_BIST_REGISTER),
    .PF1_CAPABILITY_POINTER (PF1_CAPABILITY_POINTER),
    .PF1_CLASS_CODE (PF1_CLASS_CODE),
    .PF1_DEVICE_ID (PF1_DEVICE_ID),
    .PF1_DEV_CAP_MAX_PAYLOAD_SIZE (PF1_DEV_CAP_MAX_PAYLOAD_SIZE),
    .PF1_DPA_CAP_NEXTPTR (PF1_DPA_CAP_NEXTPTR),
    .PF1_DPA_CAP_SUB_STATE_CONTROL (PF1_DPA_CAP_SUB_STATE_CONTROL),
    .PF1_DPA_CAP_SUB_STATE_CONTROL_EN (PF1_DPA_CAP_SUB_STATE_CONTROL_EN),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7),
    .PF1_DPA_CAP_VER (PF1_DPA_CAP_VER),
    .PF1_DSN_CAP_NEXTPTR (PF1_DSN_CAP_NEXTPTR),
    .PF1_EXPANSION_ROM_APERTURE_SIZE (PF1_EXPANSION_ROM_APERTURE_SIZE),
    .PF1_EXPANSION_ROM_ENABLE (PF1_EXPANSION_ROM_ENABLE),
    .PF1_INTERRUPT_LINE (PF1_INTERRUPT_LINE),
    .PF1_INTERRUPT_PIN (PF1_INTERRUPT_PIN),
    .PF1_MSIX_CAP_NEXTPTR (PF1_MSIX_CAP_NEXTPTR),
    .PF1_MSIX_CAP_PBA_BIR (PF1_MSIX_CAP_PBA_BIR),
    .PF1_MSIX_CAP_PBA_OFFSET (PF1_MSIX_CAP_PBA_OFFSET),
    .PF1_MSIX_CAP_TABLE_BIR (PF1_MSIX_CAP_TABLE_BIR),
    .PF1_MSIX_CAP_TABLE_OFFSET (PF1_MSIX_CAP_TABLE_OFFSET),
    .PF1_MSIX_CAP_TABLE_SIZE (PF1_MSIX_CAP_TABLE_SIZE),
    .PF1_MSI_CAP_MULTIMSGCAP (PF1_MSI_CAP_MULTIMSGCAP),
    .PF1_MSI_CAP_NEXTPTR (PF1_MSI_CAP_NEXTPTR),
    .PF1_PB_CAP_NEXTPTR (PF1_PB_CAP_NEXTPTR),
    .PF1_PB_CAP_SYSTEM_ALLOCATED (PF1_PB_CAP_SYSTEM_ALLOCATED),
    .PF1_PB_CAP_VER (PF1_PB_CAP_VER),
    .PF1_PM_CAP_ID (PF1_PM_CAP_ID),
    .PF1_PM_CAP_NEXTPTR (PF1_PM_CAP_NEXTPTR),
    .PF1_PM_CAP_VER_ID (PF1_PM_CAP_VER_ID),
    .PF1_RBAR_CAP_ENABLE (PF1_RBAR_CAP_ENABLE),
    .PF1_RBAR_CAP_INDEX0 (PF1_RBAR_CAP_INDEX0),
    .PF1_RBAR_CAP_INDEX1 (PF1_RBAR_CAP_INDEX1),
    .PF1_RBAR_CAP_INDEX2 (PF1_RBAR_CAP_INDEX2),
    .PF1_RBAR_CAP_NEXTPTR (PF1_RBAR_CAP_NEXTPTR),
    .PF1_RBAR_CAP_SIZE0 (PF1_RBAR_CAP_SIZE0),
    .PF1_RBAR_CAP_SIZE1 (PF1_RBAR_CAP_SIZE1),
    .PF1_RBAR_CAP_SIZE2 (PF1_RBAR_CAP_SIZE2),
    .PF1_RBAR_CAP_VER (PF1_RBAR_CAP_VER),
    .PF1_RBAR_NUM (PF1_RBAR_NUM),
    .PF1_REVISION_ID (PF1_REVISION_ID),
    .PF1_SRIOV_BAR0_APERTURE_SIZE (PF1_SRIOV_BAR0_APERTURE_SIZE),
    .PF1_SRIOV_BAR0_CONTROL (PF1_SRIOV_BAR0_CONTROL),
    .PF1_SRIOV_BAR1_APERTURE_SIZE (PF1_SRIOV_BAR1_APERTURE_SIZE),
    .PF1_SRIOV_BAR1_CONTROL (PF1_SRIOV_BAR1_CONTROL),
    .PF1_SRIOV_BAR2_APERTURE_SIZE (PF1_SRIOV_BAR2_APERTURE_SIZE),
    .PF1_SRIOV_BAR2_CONTROL (PF1_SRIOV_BAR2_CONTROL),
    .PF1_SRIOV_BAR3_APERTURE_SIZE (PF1_SRIOV_BAR3_APERTURE_SIZE),
    .PF1_SRIOV_BAR3_CONTROL (PF1_SRIOV_BAR3_CONTROL),
    .PF1_SRIOV_BAR4_APERTURE_SIZE (PF1_SRIOV_BAR4_APERTURE_SIZE),
    .PF1_SRIOV_BAR4_CONTROL (PF1_SRIOV_BAR4_CONTROL),
    .PF1_SRIOV_BAR5_APERTURE_SIZE (PF1_SRIOV_BAR5_APERTURE_SIZE),
    .PF1_SRIOV_BAR5_CONTROL (PF1_SRIOV_BAR5_CONTROL),
    .PF1_SRIOV_CAP_INITIAL_VF (PF1_SRIOV_CAP_INITIAL_VF),
    .PF1_SRIOV_CAP_NEXTPTR (PF1_SRIOV_CAP_NEXTPTR),
    .PF1_SRIOV_CAP_TOTAL_VF (PF1_SRIOV_CAP_TOTAL_VF),
    .PF1_SRIOV_CAP_VER (PF1_SRIOV_CAP_VER),
    .PF1_SRIOV_FIRST_VF_OFFSET (PF1_SRIOV_FIRST_VF_OFFSET),
    .PF1_SRIOV_FUNC_DEP_LINK (PF1_SRIOV_FUNC_DEP_LINK),
    .PF1_SRIOV_SUPPORTED_PAGE_SIZE (PF1_SRIOV_SUPPORTED_PAGE_SIZE),
    .PF1_SRIOV_VF_DEVICE_ID (PF1_SRIOV_VF_DEVICE_ID),
    .PF1_SUBSYSTEM_ID (PF1_SUBSYSTEM_ID),
    .PF1_TPHR_CAP_DEV_SPECIFIC_MODE (PF1_TPHR_CAP_DEV_SPECIFIC_MODE),
    .PF1_TPHR_CAP_ENABLE (PF1_TPHR_CAP_ENABLE),
    .PF1_TPHR_CAP_INT_VEC_MODE (PF1_TPHR_CAP_INT_VEC_MODE),
    .PF1_TPHR_CAP_NEXTPTR (PF1_TPHR_CAP_NEXTPTR),
    .PF1_TPHR_CAP_ST_MODE_SEL (PF1_TPHR_CAP_ST_MODE_SEL),
    .PF1_TPHR_CAP_ST_TABLE_LOC (PF1_TPHR_CAP_ST_TABLE_LOC),
    .PF1_TPHR_CAP_ST_TABLE_SIZE (PF1_TPHR_CAP_ST_TABLE_SIZE),
    .PF1_TPHR_CAP_VER (PF1_TPHR_CAP_VER),
    .PL_DISABLE_EI_INFER_IN_L0 (PL_DISABLE_EI_INFER_IN_L0),
    .PL_DISABLE_GEN3_DC_BALANCE (PL_DISABLE_GEN3_DC_BALANCE),
    .PL_DISABLE_SCRAMBLING (PL_DISABLE_SCRAMBLING),
    .PL_DISABLE_UPCONFIG_CAPABLE (PL_DISABLE_UPCONFIG_CAPABLE),
    .PL_EQ_ADAPT_DISABLE_COEFF_CHECK (PL_EQ_ADAPT_DISABLE_COEFF_CHECK),
    .PL_EQ_ADAPT_DISABLE_PRESET_CHECK (PL_EQ_ADAPT_DISABLE_PRESET_CHECK),
    .PL_EQ_ADAPT_ITER_COUNT (PL_EQ_ADAPT_ITER_COUNT),
    .PL_EQ_ADAPT_REJECT_RETRY_COUNT (PL_EQ_ADAPT_REJECT_RETRY_COUNT),
    .PL_EQ_BYPASS_PHASE23 (PL_EQ_BYPASS_PHASE23),
    .PL_EQ_SHORT_ADAPT_PHASE (PL_EQ_SHORT_ADAPT_PHASE),
    .PL_LANE0_EQ_CONTROL (PL_LANE0_EQ_CONTROL),
    .PL_LANE1_EQ_CONTROL (PL_LANE1_EQ_CONTROL),
    .PL_LANE2_EQ_CONTROL (PL_LANE2_EQ_CONTROL),
    .PL_LANE3_EQ_CONTROL (PL_LANE3_EQ_CONTROL),
    .PL_LANE4_EQ_CONTROL (PL_LANE4_EQ_CONTROL),
    .PL_LANE5_EQ_CONTROL (PL_LANE5_EQ_CONTROL),
    .PL_LANE6_EQ_CONTROL (PL_LANE6_EQ_CONTROL),
    .PL_LANE7_EQ_CONTROL (PL_LANE7_EQ_CONTROL),
    .PL_LINK_CAP_MAX_LINK_SPEED (PL_LINK_CAP_MAX_LINK_SPEED),
    .PL_LINK_CAP_MAX_LINK_WIDTH (PL_LINK_CAP_MAX_LINK_WIDTH),
    .PL_N_FTS_COMCLK_GEN1 (PL_N_FTS_COMCLK_GEN1),
    .PL_N_FTS_COMCLK_GEN2 (PL_N_FTS_COMCLK_GEN2),
    .PL_N_FTS_COMCLK_GEN3 (PL_N_FTS_COMCLK_GEN3),
    .PL_N_FTS_GEN1 (PL_N_FTS_GEN1),
    .PL_N_FTS_GEN2 (PL_N_FTS_GEN2),
    .PL_N_FTS_GEN3 (PL_N_FTS_GEN3),
    .PL_SIM_FAST_LINK_TRAINING (PL_SIM_FAST_LINK_TRAINING),
    .PL_UPSTREAM_FACING (PL_UPSTREAM_FACING),
    .PM_ASPML0S_TIMEOUT (PM_ASPML0S_TIMEOUT),
    .PM_ASPML1_ENTRY_DELAY (PM_ASPML1_ENTRY_DELAY),
    .PM_ENABLE_SLOT_POWER_CAPTURE (PM_ENABLE_SLOT_POWER_CAPTURE),
    .PM_L1_REENTRY_DELAY (PM_L1_REENTRY_DELAY),
    .PM_PME_SERVICE_TIMEOUT_DELAY (PM_PME_SERVICE_TIMEOUT_DELAY),
    .PM_PME_TURNOFF_ACK_DELAY (PM_PME_TURNOFF_ACK_DELAY),
    .SIM_VERSION (SIM_VERSION),
    .SPARE_BIT0 (SPARE_BIT0),
    .SPARE_BIT1 (SPARE_BIT1),
    .SPARE_BIT2 (SPARE_BIT2),
    .SPARE_BIT3 (SPARE_BIT3),
    .SPARE_BIT4 (SPARE_BIT4),
    .SPARE_BIT5 (SPARE_BIT5),
    .SPARE_BIT6 (SPARE_BIT6),
    .SPARE_BIT7 (SPARE_BIT7),
    .SPARE_BIT8 (SPARE_BIT8),
    .SPARE_BYTE0 (SPARE_BYTE0),
    .SPARE_BYTE1 (SPARE_BYTE1),
    .SPARE_BYTE2 (SPARE_BYTE2),
    .SPARE_BYTE3 (SPARE_BYTE3),
    .SPARE_WORD0 (SPARE_WORD0),
    .SPARE_WORD1 (SPARE_WORD1),
    .SPARE_WORD2 (SPARE_WORD2),
    .SPARE_WORD3 (SPARE_WORD3),
    .SRIOV_CAP_ENABLE (SRIOV_CAP_ENABLE),
    .TL_COMPL_TIMEOUT_REG0 (TL_COMPL_TIMEOUT_REG0),
    .TL_COMPL_TIMEOUT_REG1 (TL_COMPL_TIMEOUT_REG1),
    .TL_CREDITS_CD (TL_CREDITS_CD),
    .TL_CREDITS_CH (TL_CREDITS_CH),
    .TL_CREDITS_NPD (TL_CREDITS_NPD),
    .TL_CREDITS_NPH (TL_CREDITS_NPH),
    .TL_CREDITS_PD (TL_CREDITS_PD),
    .TL_CREDITS_PH (TL_CREDITS_PH),
    .TL_ENABLE_MESSAGE_RID_CHECK_ENABLE (TL_ENABLE_MESSAGE_RID_CHECK_ENABLE),
    .TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE (TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE),
    .TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE (TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE),
    .TL_LEGACY_MODE_ENABLE (TL_LEGACY_MODE_ENABLE),
    .TL_PF_ENABLE_REG (TL_PF_ENABLE_REG),
    .TL_TAG_MGMT_ENABLE (TL_TAG_MGMT_ENABLE),
    .VF0_ARI_CAP_NEXTPTR (VF0_ARI_CAP_NEXTPTR),
    .VF0_CAPABILITY_POINTER (VF0_CAPABILITY_POINTER),
    .VF0_MSIX_CAP_PBA_BIR (VF0_MSIX_CAP_PBA_BIR),
    .VF0_MSIX_CAP_PBA_OFFSET (VF0_MSIX_CAP_PBA_OFFSET),
    .VF0_MSIX_CAP_TABLE_BIR (VF0_MSIX_CAP_TABLE_BIR),
    .VF0_MSIX_CAP_TABLE_OFFSET (VF0_MSIX_CAP_TABLE_OFFSET),
    .VF0_MSIX_CAP_TABLE_SIZE (VF0_MSIX_CAP_TABLE_SIZE),
    .VF0_MSI_CAP_MULTIMSGCAP (VF0_MSI_CAP_MULTIMSGCAP),
    .VF0_PM_CAP_ID (VF0_PM_CAP_ID),
    .VF0_PM_CAP_NEXTPTR (VF0_PM_CAP_NEXTPTR),
    .VF0_PM_CAP_VER_ID (VF0_PM_CAP_VER_ID),
    .VF0_TPHR_CAP_DEV_SPECIFIC_MODE (VF0_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF0_TPHR_CAP_ENABLE (VF0_TPHR_CAP_ENABLE),
    .VF0_TPHR_CAP_INT_VEC_MODE (VF0_TPHR_CAP_INT_VEC_MODE),
    .VF0_TPHR_CAP_NEXTPTR (VF0_TPHR_CAP_NEXTPTR),
    .VF0_TPHR_CAP_ST_MODE_SEL (VF0_TPHR_CAP_ST_MODE_SEL),
    .VF0_TPHR_CAP_ST_TABLE_LOC (VF0_TPHR_CAP_ST_TABLE_LOC),
    .VF0_TPHR_CAP_ST_TABLE_SIZE (VF0_TPHR_CAP_ST_TABLE_SIZE),
    .VF0_TPHR_CAP_VER (VF0_TPHR_CAP_VER),
    .VF1_ARI_CAP_NEXTPTR (VF1_ARI_CAP_NEXTPTR),
    .VF1_MSIX_CAP_PBA_BIR (VF1_MSIX_CAP_PBA_BIR),
    .VF1_MSIX_CAP_PBA_OFFSET (VF1_MSIX_CAP_PBA_OFFSET),
    .VF1_MSIX_CAP_TABLE_BIR (VF1_MSIX_CAP_TABLE_BIR),
    .VF1_MSIX_CAP_TABLE_OFFSET (VF1_MSIX_CAP_TABLE_OFFSET),
    .VF1_MSIX_CAP_TABLE_SIZE (VF1_MSIX_CAP_TABLE_SIZE),
    .VF1_MSI_CAP_MULTIMSGCAP (VF1_MSI_CAP_MULTIMSGCAP),
    .VF1_PM_CAP_ID (VF1_PM_CAP_ID),
    .VF1_PM_CAP_NEXTPTR (VF1_PM_CAP_NEXTPTR),
    .VF1_PM_CAP_VER_ID (VF1_PM_CAP_VER_ID),
    .VF1_TPHR_CAP_DEV_SPECIFIC_MODE (VF1_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF1_TPHR_CAP_ENABLE (VF1_TPHR_CAP_ENABLE),
    .VF1_TPHR_CAP_INT_VEC_MODE (VF1_TPHR_CAP_INT_VEC_MODE),
    .VF1_TPHR_CAP_NEXTPTR (VF1_TPHR_CAP_NEXTPTR),
    .VF1_TPHR_CAP_ST_MODE_SEL (VF1_TPHR_CAP_ST_MODE_SEL),
    .VF1_TPHR_CAP_ST_TABLE_LOC (VF1_TPHR_CAP_ST_TABLE_LOC),
    .VF1_TPHR_CAP_ST_TABLE_SIZE (VF1_TPHR_CAP_ST_TABLE_SIZE),
    .VF1_TPHR_CAP_VER (VF1_TPHR_CAP_VER),
    .VF2_ARI_CAP_NEXTPTR (VF2_ARI_CAP_NEXTPTR),
    .VF2_MSIX_CAP_PBA_BIR (VF2_MSIX_CAP_PBA_BIR),
    .VF2_MSIX_CAP_PBA_OFFSET (VF2_MSIX_CAP_PBA_OFFSET),
    .VF2_MSIX_CAP_TABLE_BIR (VF2_MSIX_CAP_TABLE_BIR),
    .VF2_MSIX_CAP_TABLE_OFFSET (VF2_MSIX_CAP_TABLE_OFFSET),
    .VF2_MSIX_CAP_TABLE_SIZE (VF2_MSIX_CAP_TABLE_SIZE),
    .VF2_MSI_CAP_MULTIMSGCAP (VF2_MSI_CAP_MULTIMSGCAP),
    .VF2_PM_CAP_ID (VF2_PM_CAP_ID),
    .VF2_PM_CAP_NEXTPTR (VF2_PM_CAP_NEXTPTR),
    .VF2_PM_CAP_VER_ID (VF2_PM_CAP_VER_ID),
    .VF2_TPHR_CAP_DEV_SPECIFIC_MODE (VF2_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF2_TPHR_CAP_ENABLE (VF2_TPHR_CAP_ENABLE),
    .VF2_TPHR_CAP_INT_VEC_MODE (VF2_TPHR_CAP_INT_VEC_MODE),
    .VF2_TPHR_CAP_NEXTPTR (VF2_TPHR_CAP_NEXTPTR),
    .VF2_TPHR_CAP_ST_MODE_SEL (VF2_TPHR_CAP_ST_MODE_SEL),
    .VF2_TPHR_CAP_ST_TABLE_LOC (VF2_TPHR_CAP_ST_TABLE_LOC),
    .VF2_TPHR_CAP_ST_TABLE_SIZE (VF2_TPHR_CAP_ST_TABLE_SIZE),
    .VF2_TPHR_CAP_VER (VF2_TPHR_CAP_VER),
    .VF3_ARI_CAP_NEXTPTR (VF3_ARI_CAP_NEXTPTR),
    .VF3_MSIX_CAP_PBA_BIR (VF3_MSIX_CAP_PBA_BIR),
    .VF3_MSIX_CAP_PBA_OFFSET (VF3_MSIX_CAP_PBA_OFFSET),
    .VF3_MSIX_CAP_TABLE_BIR (VF3_MSIX_CAP_TABLE_BIR),
    .VF3_MSIX_CAP_TABLE_OFFSET (VF3_MSIX_CAP_TABLE_OFFSET),
    .VF3_MSIX_CAP_TABLE_SIZE (VF3_MSIX_CAP_TABLE_SIZE),
    .VF3_MSI_CAP_MULTIMSGCAP (VF3_MSI_CAP_MULTIMSGCAP),
    .VF3_PM_CAP_ID (VF3_PM_CAP_ID),
    .VF3_PM_CAP_NEXTPTR (VF3_PM_CAP_NEXTPTR),
    .VF3_PM_CAP_VER_ID (VF3_PM_CAP_VER_ID),
    .VF3_TPHR_CAP_DEV_SPECIFIC_MODE (VF3_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF3_TPHR_CAP_ENABLE (VF3_TPHR_CAP_ENABLE),
    .VF3_TPHR_CAP_INT_VEC_MODE (VF3_TPHR_CAP_INT_VEC_MODE),
    .VF3_TPHR_CAP_NEXTPTR (VF3_TPHR_CAP_NEXTPTR),
    .VF3_TPHR_CAP_ST_MODE_SEL (VF3_TPHR_CAP_ST_MODE_SEL),
    .VF3_TPHR_CAP_ST_TABLE_LOC (VF3_TPHR_CAP_ST_TABLE_LOC),
    .VF3_TPHR_CAP_ST_TABLE_SIZE (VF3_TPHR_CAP_ST_TABLE_SIZE),
    .VF3_TPHR_CAP_VER (VF3_TPHR_CAP_VER),
    .VF4_ARI_CAP_NEXTPTR (VF4_ARI_CAP_NEXTPTR),
    .VF4_MSIX_CAP_PBA_BIR (VF4_MSIX_CAP_PBA_BIR),
    .VF4_MSIX_CAP_PBA_OFFSET (VF4_MSIX_CAP_PBA_OFFSET),
    .VF4_MSIX_CAP_TABLE_BIR (VF4_MSIX_CAP_TABLE_BIR),
    .VF4_MSIX_CAP_TABLE_OFFSET (VF4_MSIX_CAP_TABLE_OFFSET),
    .VF4_MSIX_CAP_TABLE_SIZE (VF4_MSIX_CAP_TABLE_SIZE),
    .VF4_MSI_CAP_MULTIMSGCAP (VF4_MSI_CAP_MULTIMSGCAP),
    .VF4_PM_CAP_ID (VF4_PM_CAP_ID),
    .VF4_PM_CAP_NEXTPTR (VF4_PM_CAP_NEXTPTR),
    .VF4_PM_CAP_VER_ID (VF4_PM_CAP_VER_ID),
    .VF4_TPHR_CAP_DEV_SPECIFIC_MODE (VF4_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF4_TPHR_CAP_ENABLE (VF4_TPHR_CAP_ENABLE),
    .VF4_TPHR_CAP_INT_VEC_MODE (VF4_TPHR_CAP_INT_VEC_MODE),
    .VF4_TPHR_CAP_NEXTPTR (VF4_TPHR_CAP_NEXTPTR),
    .VF4_TPHR_CAP_ST_MODE_SEL (VF4_TPHR_CAP_ST_MODE_SEL),
    .VF4_TPHR_CAP_ST_TABLE_LOC (VF4_TPHR_CAP_ST_TABLE_LOC),
    .VF4_TPHR_CAP_ST_TABLE_SIZE (VF4_TPHR_CAP_ST_TABLE_SIZE),
    .VF4_TPHR_CAP_VER (VF4_TPHR_CAP_VER),
    .VF5_ARI_CAP_NEXTPTR (VF5_ARI_CAP_NEXTPTR),
    .VF5_MSIX_CAP_PBA_BIR (VF5_MSIX_CAP_PBA_BIR),
    .VF5_MSIX_CAP_PBA_OFFSET (VF5_MSIX_CAP_PBA_OFFSET),
    .VF5_MSIX_CAP_TABLE_BIR (VF5_MSIX_CAP_TABLE_BIR),
    .VF5_MSIX_CAP_TABLE_OFFSET (VF5_MSIX_CAP_TABLE_OFFSET),
    .VF5_MSIX_CAP_TABLE_SIZE (VF5_MSIX_CAP_TABLE_SIZE),
    .VF5_MSI_CAP_MULTIMSGCAP (VF5_MSI_CAP_MULTIMSGCAP),
    .VF5_PM_CAP_ID (VF5_PM_CAP_ID),
    .VF5_PM_CAP_NEXTPTR (VF5_PM_CAP_NEXTPTR),
    .VF5_PM_CAP_VER_ID (VF5_PM_CAP_VER_ID),
    .VF5_TPHR_CAP_DEV_SPECIFIC_MODE (VF5_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF5_TPHR_CAP_ENABLE (VF5_TPHR_CAP_ENABLE),
    .VF5_TPHR_CAP_INT_VEC_MODE (VF5_TPHR_CAP_INT_VEC_MODE),
    .VF5_TPHR_CAP_NEXTPTR (VF5_TPHR_CAP_NEXTPTR),
    .VF5_TPHR_CAP_ST_MODE_SEL (VF5_TPHR_CAP_ST_MODE_SEL),
    .VF5_TPHR_CAP_ST_TABLE_LOC (VF5_TPHR_CAP_ST_TABLE_LOC),
    .VF5_TPHR_CAP_ST_TABLE_SIZE (VF5_TPHR_CAP_ST_TABLE_SIZE),
    .VF5_TPHR_CAP_VER (VF5_TPHR_CAP_VER))

    B_PCIE_3_0_INST (
    .CFGCURRENTSPEED (delay_CFGCURRENTSPEED),
    .CFGDPASUBSTATECHANGE (delay_CFGDPASUBSTATECHANGE),
    .CFGERRCOROUT (delay_CFGERRCOROUT),
    .CFGERRFATALOUT (delay_CFGERRFATALOUT),
    .CFGERRNONFATALOUT (delay_CFGERRNONFATALOUT),
    .CFGEXTFUNCTIONNUMBER (delay_CFGEXTFUNCTIONNUMBER),
    .CFGEXTREADRECEIVED (delay_CFGEXTREADRECEIVED),
    .CFGEXTREGISTERNUMBER (delay_CFGEXTREGISTERNUMBER),
    .CFGEXTWRITEBYTEENABLE (delay_CFGEXTWRITEBYTEENABLE),
    .CFGEXTWRITEDATA (delay_CFGEXTWRITEDATA),
    .CFGEXTWRITERECEIVED (delay_CFGEXTWRITERECEIVED),
    .CFGFCCPLD (delay_CFGFCCPLD),
    .CFGFCCPLH (delay_CFGFCCPLH),
    .CFGFCNPD (delay_CFGFCNPD),
    .CFGFCNPH (delay_CFGFCNPH),
    .CFGFCPD (delay_CFGFCPD),
    .CFGFCPH (delay_CFGFCPH),
    .CFGFLRINPROCESS (delay_CFGFLRINPROCESS),
    .CFGFUNCTIONPOWERSTATE (delay_CFGFUNCTIONPOWERSTATE),
    .CFGFUNCTIONSTATUS (delay_CFGFUNCTIONSTATUS),
    .CFGHOTRESETOUT (delay_CFGHOTRESETOUT),
    .CFGINPUTUPDATEDONE (delay_CFGINPUTUPDATEDONE),
    .CFGINTERRUPTAOUTPUT (delay_CFGINTERRUPTAOUTPUT),
    .CFGINTERRUPTBOUTPUT (delay_CFGINTERRUPTBOUTPUT),
    .CFGINTERRUPTCOUTPUT (delay_CFGINTERRUPTCOUTPUT),
    .CFGINTERRUPTDOUTPUT (delay_CFGINTERRUPTDOUTPUT),
    .CFGINTERRUPTMSIDATA (delay_CFGINTERRUPTMSIDATA),
    .CFGINTERRUPTMSIENABLE (delay_CFGINTERRUPTMSIENABLE),
    .CFGINTERRUPTMSIFAIL (delay_CFGINTERRUPTMSIFAIL),
    .CFGINTERRUPTMSIMASKUPDATE (delay_CFGINTERRUPTMSIMASKUPDATE),
    .CFGINTERRUPTMSIMMENABLE (delay_CFGINTERRUPTMSIMMENABLE),
    .CFGINTERRUPTMSISENT (delay_CFGINTERRUPTMSISENT),
    .CFGINTERRUPTMSIVFENABLE (delay_CFGINTERRUPTMSIVFENABLE),
    .CFGINTERRUPTMSIXENABLE (delay_CFGINTERRUPTMSIXENABLE),
    .CFGINTERRUPTMSIXFAIL (delay_CFGINTERRUPTMSIXFAIL),
    .CFGINTERRUPTMSIXMASK (delay_CFGINTERRUPTMSIXMASK),
    .CFGINTERRUPTMSIXSENT (delay_CFGINTERRUPTMSIXSENT),
    .CFGINTERRUPTMSIXVFENABLE (delay_CFGINTERRUPTMSIXVFENABLE),
    .CFGINTERRUPTMSIXVFMASK (delay_CFGINTERRUPTMSIXVFMASK),
    .CFGINTERRUPTSENT (delay_CFGINTERRUPTSENT),
    .CFGLINKPOWERSTATE (delay_CFGLINKPOWERSTATE),
    .CFGLOCALERROR (delay_CFGLOCALERROR),
    .CFGLTRENABLE (delay_CFGLTRENABLE),
    .CFGLTSSMSTATE (delay_CFGLTSSMSTATE),
    .CFGMAXPAYLOAD (delay_CFGMAXPAYLOAD),
    .CFGMAXREADREQ (delay_CFGMAXREADREQ),
    .CFGMCUPDATEDONE (delay_CFGMCUPDATEDONE),
    .CFGMGMTREADDATA (delay_CFGMGMTREADDATA),
    .CFGMGMTREADWRITEDONE (delay_CFGMGMTREADWRITEDONE),
    .CFGMSGRECEIVED (delay_CFGMSGRECEIVED),
    .CFGMSGRECEIVEDDATA (delay_CFGMSGRECEIVEDDATA),
    .CFGMSGRECEIVEDTYPE (delay_CFGMSGRECEIVEDTYPE),
    .CFGMSGTRANSMITDONE (delay_CFGMSGTRANSMITDONE),
    .CFGNEGOTIATEDWIDTH (delay_CFGNEGOTIATEDWIDTH),
    .CFGOBFFENABLE (delay_CFGOBFFENABLE),
    .CFGPERFUNCSTATUSDATA (delay_CFGPERFUNCSTATUSDATA),
    .CFGPERFUNCTIONUPDATEDONE (delay_CFGPERFUNCTIONUPDATEDONE),
    .CFGPHYLINKDOWN (delay_CFGPHYLINKDOWN),
    .CFGPHYLINKSTATUS (delay_CFGPHYLINKSTATUS),
    .CFGPLSTATUSCHANGE (delay_CFGPLSTATUSCHANGE),
    .CFGPOWERSTATECHANGEINTERRUPT (delay_CFGPOWERSTATECHANGEINTERRUPT),
    .CFGRCBSTATUS (delay_CFGRCBSTATUS),
    .CFGTPHFUNCTIONNUM (delay_CFGTPHFUNCTIONNUM),
    .CFGTPHREQUESTERENABLE (delay_CFGTPHREQUESTERENABLE),
    .CFGTPHSTMODE (delay_CFGTPHSTMODE),
    .CFGTPHSTTADDRESS (delay_CFGTPHSTTADDRESS),
    .CFGTPHSTTREADENABLE (delay_CFGTPHSTTREADENABLE),
    .CFGTPHSTTWRITEBYTEVALID (delay_CFGTPHSTTWRITEBYTEVALID),
    .CFGTPHSTTWRITEDATA (delay_CFGTPHSTTWRITEDATA),
    .CFGTPHSTTWRITEENABLE (delay_CFGTPHSTTWRITEENABLE),
    .CFGVFFLRINPROCESS (delay_CFGVFFLRINPROCESS),
    .CFGVFPOWERSTATE (delay_CFGVFPOWERSTATE),
    .CFGVFSTATUS (delay_CFGVFSTATUS),
    .CFGVFTPHREQUESTERENABLE (delay_CFGVFTPHREQUESTERENABLE),
    .CFGVFTPHSTMODE (delay_CFGVFTPHSTMODE),
    .DBGDATAOUT (delay_DBGDATAOUT),
    .DRPDO (delay_DRPDO),
    .DRPRDY (delay_DRPRDY),
    .MAXISCQTDATA (delay_MAXISCQTDATA),
    .MAXISCQTKEEP (delay_MAXISCQTKEEP),
    .MAXISCQTLAST (delay_MAXISCQTLAST),
    .MAXISCQTUSER (delay_MAXISCQTUSER),
    .MAXISCQTVALID (delay_MAXISCQTVALID),
    .MAXISRCTDATA (delay_MAXISRCTDATA),
    .MAXISRCTKEEP (delay_MAXISRCTKEEP),
    .MAXISRCTLAST (delay_MAXISRCTLAST),
    .MAXISRCTUSER (delay_MAXISRCTUSER),
    .MAXISRCTVALID (delay_MAXISRCTVALID),
    .MICOMPLETIONRAMREADADDRESSAL (delay_MICOMPLETIONRAMREADADDRESSAL),
    .MICOMPLETIONRAMREADADDRESSAU (delay_MICOMPLETIONRAMREADADDRESSAU),
    .MICOMPLETIONRAMREADADDRESSBL (delay_MICOMPLETIONRAMREADADDRESSBL),
    .MICOMPLETIONRAMREADADDRESSBU (delay_MICOMPLETIONRAMREADADDRESSBU),
    .MICOMPLETIONRAMREADENABLEL (delay_MICOMPLETIONRAMREADENABLEL),
    .MICOMPLETIONRAMREADENABLEU (delay_MICOMPLETIONRAMREADENABLEU),
    .MICOMPLETIONRAMWRITEADDRESSAL (delay_MICOMPLETIONRAMWRITEADDRESSAL),
    .MICOMPLETIONRAMWRITEADDRESSAU (delay_MICOMPLETIONRAMWRITEADDRESSAU),
    .MICOMPLETIONRAMWRITEADDRESSBL (delay_MICOMPLETIONRAMWRITEADDRESSBL),
    .MICOMPLETIONRAMWRITEADDRESSBU (delay_MICOMPLETIONRAMWRITEADDRESSBU),
    .MICOMPLETIONRAMWRITEDATAL (delay_MICOMPLETIONRAMWRITEDATAL),
    .MICOMPLETIONRAMWRITEDATAU (delay_MICOMPLETIONRAMWRITEDATAU),
    .MICOMPLETIONRAMWRITEENABLEL (delay_MICOMPLETIONRAMWRITEENABLEL),
    .MICOMPLETIONRAMWRITEENABLEU (delay_MICOMPLETIONRAMWRITEENABLEU),
    .MIREPLAYRAMADDRESS (delay_MIREPLAYRAMADDRESS),
    .MIREPLAYRAMREADENABLE (delay_MIREPLAYRAMREADENABLE),
    .MIREPLAYRAMWRITEDATA (delay_MIREPLAYRAMWRITEDATA),
    .MIREPLAYRAMWRITEENABLE (delay_MIREPLAYRAMWRITEENABLE),
    .MIREQUESTRAMREADADDRESSA (delay_MIREQUESTRAMREADADDRESSA),
    .MIREQUESTRAMREADADDRESSB (delay_MIREQUESTRAMREADADDRESSB),
    .MIREQUESTRAMREADENABLE (delay_MIREQUESTRAMREADENABLE),
    .MIREQUESTRAMWRITEADDRESSA (delay_MIREQUESTRAMWRITEADDRESSA),
    .MIREQUESTRAMWRITEADDRESSB (delay_MIREQUESTRAMWRITEADDRESSB),
    .MIREQUESTRAMWRITEDATA (delay_MIREQUESTRAMWRITEDATA),
    .MIREQUESTRAMWRITEENABLE (delay_MIREQUESTRAMWRITEENABLE),
    .PCIECQNPREQCOUNT (delay_PCIECQNPREQCOUNT),
    .PCIERQSEQNUM (delay_PCIERQSEQNUM),
    .PCIERQSEQNUMVLD (delay_PCIERQSEQNUMVLD),
    .PCIERQTAG (delay_PCIERQTAG),
    .PCIERQTAGAV (delay_PCIERQTAGAV),
    .PCIERQTAGVLD (delay_PCIERQTAGVLD),
    .PCIETFCNPDAV (delay_PCIETFCNPDAV),
    .PCIETFCNPHAV (delay_PCIETFCNPHAV),
    .PIPERX0EQCONTROL (delay_PIPERX0EQCONTROL),
    .PIPERX0EQLPLFFS (delay_PIPERX0EQLPLFFS),
    .PIPERX0EQLPTXPRESET (delay_PIPERX0EQLPTXPRESET),
    .PIPERX0EQPRESET (delay_PIPERX0EQPRESET),
    .PIPERX0POLARITY (delay_PIPERX0POLARITY),
    .PIPERX1EQCONTROL (delay_PIPERX1EQCONTROL),
    .PIPERX1EQLPLFFS (delay_PIPERX1EQLPLFFS),
    .PIPERX1EQLPTXPRESET (delay_PIPERX1EQLPTXPRESET),
    .PIPERX1EQPRESET (delay_PIPERX1EQPRESET),
    .PIPERX1POLARITY (delay_PIPERX1POLARITY),
    .PIPERX2EQCONTROL (delay_PIPERX2EQCONTROL),
    .PIPERX2EQLPLFFS (delay_PIPERX2EQLPLFFS),
    .PIPERX2EQLPTXPRESET (delay_PIPERX2EQLPTXPRESET),
    .PIPERX2EQPRESET (delay_PIPERX2EQPRESET),
    .PIPERX2POLARITY (delay_PIPERX2POLARITY),
    .PIPERX3EQCONTROL (delay_PIPERX3EQCONTROL),
    .PIPERX3EQLPLFFS (delay_PIPERX3EQLPLFFS),
    .PIPERX3EQLPTXPRESET (delay_PIPERX3EQLPTXPRESET),
    .PIPERX3EQPRESET (delay_PIPERX3EQPRESET),
    .PIPERX3POLARITY (delay_PIPERX3POLARITY),
    .PIPERX4EQCONTROL (delay_PIPERX4EQCONTROL),
    .PIPERX4EQLPLFFS (delay_PIPERX4EQLPLFFS),
    .PIPERX4EQLPTXPRESET (delay_PIPERX4EQLPTXPRESET),
    .PIPERX4EQPRESET (delay_PIPERX4EQPRESET),
    .PIPERX4POLARITY (delay_PIPERX4POLARITY),
    .PIPERX5EQCONTROL (delay_PIPERX5EQCONTROL),
    .PIPERX5EQLPLFFS (delay_PIPERX5EQLPLFFS),
    .PIPERX5EQLPTXPRESET (delay_PIPERX5EQLPTXPRESET),
    .PIPERX5EQPRESET (delay_PIPERX5EQPRESET),
    .PIPERX5POLARITY (delay_PIPERX5POLARITY),
    .PIPERX6EQCONTROL (delay_PIPERX6EQCONTROL),
    .PIPERX6EQLPLFFS (delay_PIPERX6EQLPLFFS),
    .PIPERX6EQLPTXPRESET (delay_PIPERX6EQLPTXPRESET),
    .PIPERX6EQPRESET (delay_PIPERX6EQPRESET),
    .PIPERX6POLARITY (delay_PIPERX6POLARITY),
    .PIPERX7EQCONTROL (delay_PIPERX7EQCONTROL),
    .PIPERX7EQLPLFFS (delay_PIPERX7EQLPLFFS),
    .PIPERX7EQLPTXPRESET (delay_PIPERX7EQLPTXPRESET),
    .PIPERX7EQPRESET (delay_PIPERX7EQPRESET),
    .PIPERX7POLARITY (delay_PIPERX7POLARITY),
    .PIPETX0CHARISK (delay_PIPETX0CHARISK),
    .PIPETX0COMPLIANCE (delay_PIPETX0COMPLIANCE),
    .PIPETX0DATA (delay_PIPETX0DATA),
    .PIPETX0DATAVALID (delay_PIPETX0DATAVALID),
    .PIPETX0ELECIDLE (delay_PIPETX0ELECIDLE),
    .PIPETX0EQCONTROL (delay_PIPETX0EQCONTROL),
    .PIPETX0EQDEEMPH (delay_PIPETX0EQDEEMPH),
    .PIPETX0EQPRESET (delay_PIPETX0EQPRESET),
    .PIPETX0POWERDOWN (delay_PIPETX0POWERDOWN),
    .PIPETX0STARTBLOCK (delay_PIPETX0STARTBLOCK),
    .PIPETX0SYNCHEADER (delay_PIPETX0SYNCHEADER),
    .PIPETX1CHARISK (delay_PIPETX1CHARISK),
    .PIPETX1COMPLIANCE (delay_PIPETX1COMPLIANCE),
    .PIPETX1DATA (delay_PIPETX1DATA),
    .PIPETX1DATAVALID (delay_PIPETX1DATAVALID),
    .PIPETX1ELECIDLE (delay_PIPETX1ELECIDLE),
    .PIPETX1EQCONTROL (delay_PIPETX1EQCONTROL),
    .PIPETX1EQDEEMPH (delay_PIPETX1EQDEEMPH),
    .PIPETX1EQPRESET (delay_PIPETX1EQPRESET),
    .PIPETX1POWERDOWN (delay_PIPETX1POWERDOWN),
    .PIPETX1STARTBLOCK (delay_PIPETX1STARTBLOCK),
    .PIPETX1SYNCHEADER (delay_PIPETX1SYNCHEADER),
    .PIPETX2CHARISK (delay_PIPETX2CHARISK),
    .PIPETX2COMPLIANCE (delay_PIPETX2COMPLIANCE),
    .PIPETX2DATA (delay_PIPETX2DATA),
    .PIPETX2DATAVALID (delay_PIPETX2DATAVALID),
    .PIPETX2ELECIDLE (delay_PIPETX2ELECIDLE),
    .PIPETX2EQCONTROL (delay_PIPETX2EQCONTROL),
    .PIPETX2EQDEEMPH (delay_PIPETX2EQDEEMPH),
    .PIPETX2EQPRESET (delay_PIPETX2EQPRESET),
    .PIPETX2POWERDOWN (delay_PIPETX2POWERDOWN),
    .PIPETX2STARTBLOCK (delay_PIPETX2STARTBLOCK),
    .PIPETX2SYNCHEADER (delay_PIPETX2SYNCHEADER),
    .PIPETX3CHARISK (delay_PIPETX3CHARISK),
    .PIPETX3COMPLIANCE (delay_PIPETX3COMPLIANCE),
    .PIPETX3DATA (delay_PIPETX3DATA),
    .PIPETX3DATAVALID (delay_PIPETX3DATAVALID),
    .PIPETX3ELECIDLE (delay_PIPETX3ELECIDLE),
    .PIPETX3EQCONTROL (delay_PIPETX3EQCONTROL),
    .PIPETX3EQDEEMPH (delay_PIPETX3EQDEEMPH),
    .PIPETX3EQPRESET (delay_PIPETX3EQPRESET),
    .PIPETX3POWERDOWN (delay_PIPETX3POWERDOWN),
    .PIPETX3STARTBLOCK (delay_PIPETX3STARTBLOCK),
    .PIPETX3SYNCHEADER (delay_PIPETX3SYNCHEADER),
    .PIPETX4CHARISK (delay_PIPETX4CHARISK),
    .PIPETX4COMPLIANCE (delay_PIPETX4COMPLIANCE),
    .PIPETX4DATA (delay_PIPETX4DATA),
    .PIPETX4DATAVALID (delay_PIPETX4DATAVALID),
    .PIPETX4ELECIDLE (delay_PIPETX4ELECIDLE),
    .PIPETX4EQCONTROL (delay_PIPETX4EQCONTROL),
    .PIPETX4EQDEEMPH (delay_PIPETX4EQDEEMPH),
    .PIPETX4EQPRESET (delay_PIPETX4EQPRESET),
    .PIPETX4POWERDOWN (delay_PIPETX4POWERDOWN),
    .PIPETX4STARTBLOCK (delay_PIPETX4STARTBLOCK),
    .PIPETX4SYNCHEADER (delay_PIPETX4SYNCHEADER),
    .PIPETX5CHARISK (delay_PIPETX5CHARISK),
    .PIPETX5COMPLIANCE (delay_PIPETX5COMPLIANCE),
    .PIPETX5DATA (delay_PIPETX5DATA),
    .PIPETX5DATAVALID (delay_PIPETX5DATAVALID),
    .PIPETX5ELECIDLE (delay_PIPETX5ELECIDLE),
    .PIPETX5EQCONTROL (delay_PIPETX5EQCONTROL),
    .PIPETX5EQDEEMPH (delay_PIPETX5EQDEEMPH),
    .PIPETX5EQPRESET (delay_PIPETX5EQPRESET),
    .PIPETX5POWERDOWN (delay_PIPETX5POWERDOWN),
    .PIPETX5STARTBLOCK (delay_PIPETX5STARTBLOCK),
    .PIPETX5SYNCHEADER (delay_PIPETX5SYNCHEADER),
    .PIPETX6CHARISK (delay_PIPETX6CHARISK),
    .PIPETX6COMPLIANCE (delay_PIPETX6COMPLIANCE),
    .PIPETX6DATA (delay_PIPETX6DATA),
    .PIPETX6DATAVALID (delay_PIPETX6DATAVALID),
    .PIPETX6ELECIDLE (delay_PIPETX6ELECIDLE),
    .PIPETX6EQCONTROL (delay_PIPETX6EQCONTROL),
    .PIPETX6EQDEEMPH (delay_PIPETX6EQDEEMPH),
    .PIPETX6EQPRESET (delay_PIPETX6EQPRESET),
    .PIPETX6POWERDOWN (delay_PIPETX6POWERDOWN),
    .PIPETX6STARTBLOCK (delay_PIPETX6STARTBLOCK),
    .PIPETX6SYNCHEADER (delay_PIPETX6SYNCHEADER),
    .PIPETX7CHARISK (delay_PIPETX7CHARISK),
    .PIPETX7COMPLIANCE (delay_PIPETX7COMPLIANCE),
    .PIPETX7DATA (delay_PIPETX7DATA),
    .PIPETX7DATAVALID (delay_PIPETX7DATAVALID),
    .PIPETX7ELECIDLE (delay_PIPETX7ELECIDLE),
    .PIPETX7EQCONTROL (delay_PIPETX7EQCONTROL),
    .PIPETX7EQDEEMPH (delay_PIPETX7EQDEEMPH),
    .PIPETX7EQPRESET (delay_PIPETX7EQPRESET),
    .PIPETX7POWERDOWN (delay_PIPETX7POWERDOWN),
    .PIPETX7STARTBLOCK (delay_PIPETX7STARTBLOCK),
    .PIPETX7SYNCHEADER (delay_PIPETX7SYNCHEADER),
    .PIPETXDEEMPH (delay_PIPETXDEEMPH),
    .PIPETXMARGIN (delay_PIPETXMARGIN),
    .PIPETXRATE (delay_PIPETXRATE),
    .PIPETXRCVRDET (delay_PIPETXRCVRDET),
    .PIPETXRESET (delay_PIPETXRESET),
    .PIPETXSWING (delay_PIPETXSWING),
    .PLEQINPROGRESS (delay_PLEQINPROGRESS),
    .PLEQPHASE (delay_PLEQPHASE),
    .PLGEN3PCSRXSLIDE (delay_PLGEN3PCSRXSLIDE),
    .SAXISCCTREADY (delay_SAXISCCTREADY),
    .SAXISRQTREADY (delay_SAXISRQTREADY),
    .CFGCONFIGSPACEENABLE (delay_CFGCONFIGSPACEENABLE),
    .CFGDEVID (delay_CFGDEVID),
    .CFGDSBUSNUMBER (delay_CFGDSBUSNUMBER),
    .CFGDSDEVICENUMBER (delay_CFGDSDEVICENUMBER),
    .CFGDSFUNCTIONNUMBER (delay_CFGDSFUNCTIONNUMBER),
    .CFGDSN (delay_CFGDSN),
    .CFGDSPORTNUMBER (delay_CFGDSPORTNUMBER),
    .CFGERRCORIN (delay_CFGERRCORIN),
    .CFGERRUNCORIN (delay_CFGERRUNCORIN),
    .CFGEXTREADDATA (delay_CFGEXTREADDATA),
    .CFGEXTREADDATAVALID (delay_CFGEXTREADDATAVALID),
    .CFGFCSEL (delay_CFGFCSEL),
    .CFGFLRDONE (delay_CFGFLRDONE),
    .CFGHOTRESETIN (delay_CFGHOTRESETIN),
    .CFGINPUTUPDATEREQUEST (delay_CFGINPUTUPDATEREQUEST),
    .CFGINTERRUPTINT (delay_CFGINTERRUPTINT),
    .CFGINTERRUPTMSIATTR (delay_CFGINTERRUPTMSIATTR),
    .CFGINTERRUPTMSIFUNCTIONNUMBER (delay_CFGINTERRUPTMSIFUNCTIONNUMBER),
    .CFGINTERRUPTMSIINT (delay_CFGINTERRUPTMSIINT),
    .CFGINTERRUPTMSIPENDINGSTATUS (delay_CFGINTERRUPTMSIPENDINGSTATUS),
    .CFGINTERRUPTMSISELECT (delay_CFGINTERRUPTMSISELECT),
    .CFGINTERRUPTMSITPHPRESENT (delay_CFGINTERRUPTMSITPHPRESENT),
    .CFGINTERRUPTMSITPHSTTAG (delay_CFGINTERRUPTMSITPHSTTAG),
    .CFGINTERRUPTMSITPHTYPE (delay_CFGINTERRUPTMSITPHTYPE),
    .CFGINTERRUPTMSIXADDRESS (delay_CFGINTERRUPTMSIXADDRESS),
    .CFGINTERRUPTMSIXDATA (delay_CFGINTERRUPTMSIXDATA),
    .CFGINTERRUPTMSIXINT (delay_CFGINTERRUPTMSIXINT),
    .CFGINTERRUPTPENDING (delay_CFGINTERRUPTPENDING),
    .CFGLINKTRAININGENABLE (delay_CFGLINKTRAININGENABLE),
    .CFGMCUPDATEREQUEST (delay_CFGMCUPDATEREQUEST),
    .CFGMGMTADDR (delay_CFGMGMTADDR),
    .CFGMGMTBYTEENABLE (delay_CFGMGMTBYTEENABLE),
    .CFGMGMTREAD (delay_CFGMGMTREAD),
    .CFGMGMTTYPE1CFGREGACCESS (delay_CFGMGMTTYPE1CFGREGACCESS),
    .CFGMGMTWRITE (delay_CFGMGMTWRITE),
    .CFGMGMTWRITEDATA (delay_CFGMGMTWRITEDATA),
    .CFGMSGTRANSMIT (delay_CFGMSGTRANSMIT),
    .CFGMSGTRANSMITDATA (delay_CFGMSGTRANSMITDATA),
    .CFGMSGTRANSMITTYPE (delay_CFGMSGTRANSMITTYPE),
    .CFGPERFUNCSTATUSCONTROL (delay_CFGPERFUNCSTATUSCONTROL),
    .CFGPERFUNCTIONNUMBER (delay_CFGPERFUNCTIONNUMBER),
    .CFGPERFUNCTIONOUTPUTREQUEST (delay_CFGPERFUNCTIONOUTPUTREQUEST),
    .CFGPOWERSTATECHANGEACK (delay_CFGPOWERSTATECHANGEACK),
    .CFGREQPMTRANSITIONL23READY (delay_CFGREQPMTRANSITIONL23READY),
    .CFGREVID (delay_CFGREVID),
    .CFGSUBSYSID (delay_CFGSUBSYSID),
    .CFGSUBSYSVENDID (delay_CFGSUBSYSVENDID),
    .CFGTPHSTTREADDATA (delay_CFGTPHSTTREADDATA),
    .CFGTPHSTTREADDATAVALID (delay_CFGTPHSTTREADDATAVALID),
    .CFGVENDID (delay_CFGVENDID),
    .CFGVFFLRDONE (delay_CFGVFFLRDONE),
    .CORECLK (delay_CORECLK),
    .CORECLKMICOMPLETIONRAML (delay_CORECLKMICOMPLETIONRAML),
    .CORECLKMICOMPLETIONRAMU (delay_CORECLKMICOMPLETIONRAMU),
    .CORECLKMIREPLAYRAM (delay_CORECLKMIREPLAYRAM),
    .CORECLKMIREQUESTRAM (delay_CORECLKMIREQUESTRAM),
    .DRPADDR (delay_DRPADDR),
    .DRPCLK (delay_DRPCLK),
    .DRPDI (delay_DRPDI),
    .DRPEN (delay_DRPEN),
    .DRPWE (delay_DRPWE),
    .MAXISCQTREADY (delay_MAXISCQTREADY),
    .MAXISRCTREADY (delay_MAXISRCTREADY),
    .MGMTRESETN (delay_MGMTRESETN),
    .MGMTSTICKYRESETN (delay_MGMTSTICKYRESETN),
    .MICOMPLETIONRAMREADDATA (delay_MICOMPLETIONRAMREADDATA),
    .MIREPLAYRAMREADDATA (delay_MIREPLAYRAMREADDATA),
    .MIREQUESTRAMREADDATA (delay_MIREQUESTRAMREADDATA),
    .PCIECQNPREQ (delay_PCIECQNPREQ),
    .PIPECLK (delay_PIPECLK),
    .PIPEEQFS (delay_PIPEEQFS),
    .PIPEEQLF (delay_PIPEEQLF),
    .PIPERESETN (delay_PIPERESETN),
    .PIPERX0CHARISK (delay_PIPERX0CHARISK),
    .PIPERX0DATA (delay_PIPERX0DATA),
    .PIPERX0DATAVALID (delay_PIPERX0DATAVALID),
    .PIPERX0ELECIDLE (delay_PIPERX0ELECIDLE),
    .PIPERX0EQDONE (delay_PIPERX0EQDONE),
    .PIPERX0EQLPADAPTDONE (delay_PIPERX0EQLPADAPTDONE),
    .PIPERX0EQLPLFFSSEL (delay_PIPERX0EQLPLFFSSEL),
    .PIPERX0EQLPNEWTXCOEFFORPRESET (delay_PIPERX0EQLPNEWTXCOEFFORPRESET),
    .PIPERX0PHYSTATUS (delay_PIPERX0PHYSTATUS),
    .PIPERX0STARTBLOCK (delay_PIPERX0STARTBLOCK),
    .PIPERX0STATUS (delay_PIPERX0STATUS),
    .PIPERX0SYNCHEADER (delay_PIPERX0SYNCHEADER),
    .PIPERX0VALID (delay_PIPERX0VALID),
    .PIPERX1CHARISK (delay_PIPERX1CHARISK),
    .PIPERX1DATA (delay_PIPERX1DATA),
    .PIPERX1DATAVALID (delay_PIPERX1DATAVALID),
    .PIPERX1ELECIDLE (delay_PIPERX1ELECIDLE),
    .PIPERX1EQDONE (delay_PIPERX1EQDONE),
    .PIPERX1EQLPADAPTDONE (delay_PIPERX1EQLPADAPTDONE),
    .PIPERX1EQLPLFFSSEL (delay_PIPERX1EQLPLFFSSEL),
    .PIPERX1EQLPNEWTXCOEFFORPRESET (delay_PIPERX1EQLPNEWTXCOEFFORPRESET),
    .PIPERX1PHYSTATUS (delay_PIPERX1PHYSTATUS),
    .PIPERX1STARTBLOCK (delay_PIPERX1STARTBLOCK),
    .PIPERX1STATUS (delay_PIPERX1STATUS),
    .PIPERX1SYNCHEADER (delay_PIPERX1SYNCHEADER),
    .PIPERX1VALID (delay_PIPERX1VALID),
    .PIPERX2CHARISK (delay_PIPERX2CHARISK),
    .PIPERX2DATA (delay_PIPERX2DATA),
    .PIPERX2DATAVALID (delay_PIPERX2DATAVALID),
    .PIPERX2ELECIDLE (delay_PIPERX2ELECIDLE),
    .PIPERX2EQDONE (delay_PIPERX2EQDONE),
    .PIPERX2EQLPADAPTDONE (delay_PIPERX2EQLPADAPTDONE),
    .PIPERX2EQLPLFFSSEL (delay_PIPERX2EQLPLFFSSEL),
    .PIPERX2EQLPNEWTXCOEFFORPRESET (delay_PIPERX2EQLPNEWTXCOEFFORPRESET),
    .PIPERX2PHYSTATUS (delay_PIPERX2PHYSTATUS),
    .PIPERX2STARTBLOCK (delay_PIPERX2STARTBLOCK),
    .PIPERX2STATUS (delay_PIPERX2STATUS),
    .PIPERX2SYNCHEADER (delay_PIPERX2SYNCHEADER),
    .PIPERX2VALID (delay_PIPERX2VALID),
    .PIPERX3CHARISK (delay_PIPERX3CHARISK),
    .PIPERX3DATA (delay_PIPERX3DATA),
    .PIPERX3DATAVALID (delay_PIPERX3DATAVALID),
    .PIPERX3ELECIDLE (delay_PIPERX3ELECIDLE),
    .PIPERX3EQDONE (delay_PIPERX3EQDONE),
    .PIPERX3EQLPADAPTDONE (delay_PIPERX3EQLPADAPTDONE),
    .PIPERX3EQLPLFFSSEL (delay_PIPERX3EQLPLFFSSEL),
    .PIPERX3EQLPNEWTXCOEFFORPRESET (delay_PIPERX3EQLPNEWTXCOEFFORPRESET),
    .PIPERX3PHYSTATUS (delay_PIPERX3PHYSTATUS),
    .PIPERX3STARTBLOCK (delay_PIPERX3STARTBLOCK),
    .PIPERX3STATUS (delay_PIPERX3STATUS),
    .PIPERX3SYNCHEADER (delay_PIPERX3SYNCHEADER),
    .PIPERX3VALID (delay_PIPERX3VALID),
    .PIPERX4CHARISK (delay_PIPERX4CHARISK),
    .PIPERX4DATA (delay_PIPERX4DATA),
    .PIPERX4DATAVALID (delay_PIPERX4DATAVALID),
    .PIPERX4ELECIDLE (delay_PIPERX4ELECIDLE),
    .PIPERX4EQDONE (delay_PIPERX4EQDONE),
    .PIPERX4EQLPADAPTDONE (delay_PIPERX4EQLPADAPTDONE),
    .PIPERX4EQLPLFFSSEL (delay_PIPERX4EQLPLFFSSEL),
    .PIPERX4EQLPNEWTXCOEFFORPRESET (delay_PIPERX4EQLPNEWTXCOEFFORPRESET),
    .PIPERX4PHYSTATUS (delay_PIPERX4PHYSTATUS),
    .PIPERX4STARTBLOCK (delay_PIPERX4STARTBLOCK),
    .PIPERX4STATUS (delay_PIPERX4STATUS),
    .PIPERX4SYNCHEADER (delay_PIPERX4SYNCHEADER),
    .PIPERX4VALID (delay_PIPERX4VALID),
    .PIPERX5CHARISK (delay_PIPERX5CHARISK),
    .PIPERX5DATA (delay_PIPERX5DATA),
    .PIPERX5DATAVALID (delay_PIPERX5DATAVALID),
    .PIPERX5ELECIDLE (delay_PIPERX5ELECIDLE),
    .PIPERX5EQDONE (delay_PIPERX5EQDONE),
    .PIPERX5EQLPADAPTDONE (delay_PIPERX5EQLPADAPTDONE),
    .PIPERX5EQLPLFFSSEL (delay_PIPERX5EQLPLFFSSEL),
    .PIPERX5EQLPNEWTXCOEFFORPRESET (delay_PIPERX5EQLPNEWTXCOEFFORPRESET),
    .PIPERX5PHYSTATUS (delay_PIPERX5PHYSTATUS),
    .PIPERX5STARTBLOCK (delay_PIPERX5STARTBLOCK),
    .PIPERX5STATUS (delay_PIPERX5STATUS),
    .PIPERX5SYNCHEADER (delay_PIPERX5SYNCHEADER),
    .PIPERX5VALID (delay_PIPERX5VALID),
    .PIPERX6CHARISK (delay_PIPERX6CHARISK),
    .PIPERX6DATA (delay_PIPERX6DATA),
    .PIPERX6DATAVALID (delay_PIPERX6DATAVALID),
    .PIPERX6ELECIDLE (delay_PIPERX6ELECIDLE),
    .PIPERX6EQDONE (delay_PIPERX6EQDONE),
    .PIPERX6EQLPADAPTDONE (delay_PIPERX6EQLPADAPTDONE),
    .PIPERX6EQLPLFFSSEL (delay_PIPERX6EQLPLFFSSEL),
    .PIPERX6EQLPNEWTXCOEFFORPRESET (delay_PIPERX6EQLPNEWTXCOEFFORPRESET),
    .PIPERX6PHYSTATUS (delay_PIPERX6PHYSTATUS),
    .PIPERX6STARTBLOCK (delay_PIPERX6STARTBLOCK),
    .PIPERX6STATUS (delay_PIPERX6STATUS),
    .PIPERX6SYNCHEADER (delay_PIPERX6SYNCHEADER),
    .PIPERX6VALID (delay_PIPERX6VALID),
    .PIPERX7CHARISK (delay_PIPERX7CHARISK),
    .PIPERX7DATA (delay_PIPERX7DATA),
    .PIPERX7DATAVALID (delay_PIPERX7DATAVALID),
    .PIPERX7ELECIDLE (delay_PIPERX7ELECIDLE),
    .PIPERX7EQDONE (delay_PIPERX7EQDONE),
    .PIPERX7EQLPADAPTDONE (delay_PIPERX7EQLPADAPTDONE),
    .PIPERX7EQLPLFFSSEL (delay_PIPERX7EQLPLFFSSEL),
    .PIPERX7EQLPNEWTXCOEFFORPRESET (delay_PIPERX7EQLPNEWTXCOEFFORPRESET),
    .PIPERX7PHYSTATUS (delay_PIPERX7PHYSTATUS),
    .PIPERX7STARTBLOCK (delay_PIPERX7STARTBLOCK),
    .PIPERX7STATUS (delay_PIPERX7STATUS),
    .PIPERX7SYNCHEADER (delay_PIPERX7SYNCHEADER),
    .PIPERX7VALID (delay_PIPERX7VALID),
    .PIPETX0EQCOEFF (delay_PIPETX0EQCOEFF),
    .PIPETX0EQDONE (delay_PIPETX0EQDONE),
    .PIPETX1EQCOEFF (delay_PIPETX1EQCOEFF),
    .PIPETX1EQDONE (delay_PIPETX1EQDONE),
    .PIPETX2EQCOEFF (delay_PIPETX2EQCOEFF),
    .PIPETX2EQDONE (delay_PIPETX2EQDONE),
    .PIPETX3EQCOEFF (delay_PIPETX3EQCOEFF),
    .PIPETX3EQDONE (delay_PIPETX3EQDONE),
    .PIPETX4EQCOEFF (delay_PIPETX4EQCOEFF),
    .PIPETX4EQDONE (delay_PIPETX4EQDONE),
    .PIPETX5EQCOEFF (delay_PIPETX5EQCOEFF),
    .PIPETX5EQDONE (delay_PIPETX5EQDONE),
    .PIPETX6EQCOEFF (delay_PIPETX6EQCOEFF),
    .PIPETX6EQDONE (delay_PIPETX6EQDONE),
    .PIPETX7EQCOEFF (delay_PIPETX7EQCOEFF),
    .PIPETX7EQDONE (delay_PIPETX7EQDONE),
    .PLDISABLESCRAMBLER (delay_PLDISABLESCRAMBLER),
    .PLEQRESETEIEOSCOUNT (delay_PLEQRESETEIEOSCOUNT),
    .PLGEN3PCSDISABLE (delay_PLGEN3PCSDISABLE),
    .PLGEN3PCSRXSYNCDONE (delay_PLGEN3PCSRXSYNCDONE),
    .RECCLK (delay_RECCLK),
    .RESETN (delay_RESETN),
    .SAXISCCTDATA (delay_SAXISCCTDATA),
    .SAXISCCTKEEP (delay_SAXISCCTKEEP),
    .SAXISCCTLAST (delay_SAXISCCTLAST),
    .SAXISCCTUSER (delay_SAXISCCTUSER),
    .SAXISCCTVALID (delay_SAXISCCTVALID),
    .SAXISRQTDATA (delay_SAXISRQTDATA),
    .SAXISRQTKEEP (delay_SAXISRQTKEEP),
    .SAXISRQTLAST (delay_SAXISRQTLAST),
    .SAXISRQTUSER (delay_SAXISRQTUSER),
    .SAXISRQTVALID (delay_SAXISRQTVALID),
    .USERCLK (delay_USERCLK)
  );

  specify
`ifdef XIL_TIMING // Simprim
    $period (posedge CORECLK, 0:0:0, notifier);
    $period (posedge CORECLKMICOMPLETIONRAML, 0:0:0, notifier);
    $period (posedge CORECLKMICOMPLETIONRAMU, 0:0:0, notifier);
    $period (posedge CORECLKMIREPLAYRAM, 0:0:0, notifier);
    $period (posedge CORECLKMIREQUESTRAM, 0:0:0, notifier);
    $period (posedge DRPCLK, 0:0:0, notifier);
    $period (posedge PIPECLK, 0:0:0, notifier);
    $period (posedge RECCLK, 0:0:0, notifier);
    $period (posedge USERCLK, 0:0:0, notifier);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[0]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[100]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[101]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[102]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[103]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[104]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[105]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[106]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[107]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[108]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[109]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[10]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[110]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[111]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[112]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[113]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[114]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[115]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[116]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[117]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[118]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[119]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[11]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[120]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[121]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[122]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[123]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[124]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[125]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[126]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[127]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[128]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[129]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[12]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[130]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[131]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[132]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[133]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[134]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[135]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[136]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[137]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[138]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[139]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[13]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[140]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[141]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[142]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[143]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[14]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[15]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[16]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[17]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[18]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[19]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[1]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[20]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[21]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[22]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[23]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[24]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[25]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[26]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[27]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[28]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[29]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[2]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[30]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[31]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[32]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[33]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[34]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[35]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[36]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[37]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[38]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[39]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[3]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[40]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[41]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[42]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[43]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[44]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[45]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[46]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[47]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[48]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[49]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[4]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[50]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[51]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[52]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[53]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[54]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[55]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[56]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[57]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[58]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[59]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[5]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[60]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[61]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[62]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[63]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[64]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[65]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[66]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[67]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[68]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[69]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[6]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[70]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[71]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[72]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[73]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[74]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[75]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[76]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[77]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[78]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[79]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[7]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[80]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[81]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[82]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[83]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[84]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[85]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[86]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[87]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[88]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[89]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[8]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[90]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[91]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[92]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[93]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[94]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[95]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[96]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[97]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[98]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[99]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[9]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[0]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[100]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[101]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[102]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[103]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[104]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[105]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[106]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[107]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[108]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[109]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[10]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[110]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[111]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[112]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[113]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[114]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[115]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[116]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[117]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[118]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[119]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[11]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[120]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[121]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[122]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[123]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[124]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[125]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[126]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[127]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[128]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[129]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[12]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[130]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[131]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[132]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[133]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[134]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[135]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[136]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[137]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[138]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[139]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[13]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[140]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[141]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[142]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[143]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[14]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[15]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[16]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[17]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[18]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[19]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[1]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[20]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[21]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[22]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[23]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[24]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[25]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[26]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[27]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[28]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[29]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[2]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[30]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[31]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[32]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[33]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[34]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[35]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[36]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[37]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[38]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[39]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[3]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[40]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[41]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[42]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[43]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[44]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[45]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[46]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[47]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[48]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[49]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[4]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[50]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[51]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[52]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[53]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[54]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[55]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[56]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[57]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[58]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[59]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[5]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[60]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[61]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[62]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[63]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[64]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[65]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[66]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[67]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[68]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[69]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[6]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[70]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[71]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[72]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[73]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[74]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[75]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[76]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[77]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[78]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[79]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[7]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[80]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[81]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[82]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[83]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[84]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[85]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[86]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[87]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[88]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[89]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[8]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[90]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[91]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[92]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[93]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[94]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[95]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[96]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[97]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[98]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[99]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[9]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[0]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[100]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[101]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[102]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[103]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[104]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[105]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[106]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[107]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[108]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[109]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[10]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[110]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[111]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[112]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[113]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[114]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[115]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[116]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[117]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[118]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[119]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[11]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[120]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[121]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[122]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[123]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[124]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[125]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[126]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[127]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[128]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[129]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[12]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[130]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[131]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[132]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[133]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[134]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[135]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[136]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[137]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[138]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[139]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[13]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[140]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[141]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[142]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[143]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[14]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[15]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[16]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[17]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[18]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[19]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[1]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[20]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[21]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[22]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[23]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[24]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[25]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[26]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[27]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[28]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[29]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[2]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[30]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[31]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[32]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[33]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[34]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[35]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[36]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[37]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[38]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[39]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[3]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[40]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[41]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[42]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[43]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[44]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[45]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[46]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[47]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[48]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[49]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[4]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[50]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[51]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[52]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[53]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[54]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[55]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[56]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[57]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[58]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[59]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[5]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[60]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[61]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[62]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[63]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[64]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[65]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[66]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[67]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[68]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[69]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[6]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[70]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[71]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[72]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[73]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[74]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[75]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[76]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[77]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[78]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[79]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[7]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[80]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[81]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[82]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[83]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[84]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[85]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[86]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[87]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[88]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[89]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[8]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[90]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[91]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[92]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[93]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[94]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[95]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[96]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[97]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[98]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[99]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[9]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[0]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[100]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[101]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[102]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[103]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[104]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[105]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[106]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[107]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[108]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[109]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[10]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[110]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[111]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[112]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[113]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[114]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[115]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[116]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[117]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[118]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[119]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[11]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[120]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[121]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[122]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[123]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[124]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[125]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[126]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[127]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[128]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[129]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[12]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[130]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[131]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[132]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[133]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[134]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[135]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[136]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[137]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[138]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[139]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[13]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[140]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[141]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[142]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[143]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[14]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[15]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[16]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[17]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[18]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[19]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[1]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[20]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[21]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[22]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[23]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[24]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[25]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[26]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[27]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[28]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[29]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[2]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[30]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[31]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[32]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[33]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[34]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[35]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[36]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[37]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[38]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[39]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[3]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[40]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[41]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[42]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[43]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[44]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[45]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[46]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[47]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[48]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[49]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[4]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[50]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[51]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[52]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[53]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[54]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[55]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[56]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[57]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[58]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[59]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[5]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[60]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[61]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[62]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[63]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[64]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[65]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[66]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[67]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[68]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[69]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[6]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[70]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[71]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[72]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[73]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[74]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[75]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[76]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[77]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[78]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[79]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[7]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[80]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[81]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[82]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[83]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[84]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[85]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[86]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[87]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[88]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[89]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[8]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[90]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[91]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[92]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[93]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[94]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[95]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[96]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[97]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[98]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[99]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[9]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[0]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[100]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[101]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[102]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[103]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[104]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[105]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[106]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[107]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[108]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[109]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[10]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[110]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[111]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[112]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[113]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[114]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[115]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[116]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[117]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[118]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[119]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[11]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[120]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[121]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[122]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[123]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[124]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[125]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[126]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[127]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[128]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[129]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[12]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[130]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[131]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[132]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[133]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[134]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[135]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[136]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[137]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[138]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[139]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[13]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[140]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[141]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[142]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[143]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[14]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[15]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[16]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[17]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[18]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[19]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[1]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[20]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[21]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[22]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[23]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[24]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[25]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[26]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[27]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[28]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[29]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[2]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[30]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[31]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[32]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[33]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[34]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[35]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[36]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[37]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[38]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[39]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[3]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[40]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[41]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[42]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[43]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[44]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[45]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[46]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[47]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[48]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[49]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[4]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[50]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[51]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[52]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[53]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[54]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[55]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[56]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[57]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[58]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[59]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[5]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[60]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[61]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[62]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[63]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[64]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[65]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[66]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[67]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[68]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[69]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[6]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[70]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[71]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[72]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[73]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[74]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[75]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[76]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[77]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[78]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[79]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[7]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[80]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[81]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[82]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[83]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[84]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[85]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[86]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[87]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[88]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[89]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[8]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[90]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[91]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[92]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[93]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[94]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[95]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[96]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[97]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[98]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[99]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[9]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[0]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[100]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[101]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[102]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[103]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[104]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[105]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[106]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[107]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[108]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[109]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[10]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[110]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[111]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[112]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[113]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[114]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[115]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[116]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[117]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[118]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[119]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[11]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[120]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[121]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[122]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[123]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[124]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[125]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[126]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[127]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[128]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[129]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[12]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[130]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[131]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[132]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[133]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[134]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[135]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[136]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[137]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[138]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[139]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[13]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[140]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[141]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[142]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[143]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[14]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[15]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[16]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[17]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[18]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[19]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[1]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[20]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[21]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[22]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[23]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[24]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[25]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[26]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[27]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[28]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[29]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[2]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[30]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[31]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[32]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[33]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[34]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[35]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[36]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[37]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[38]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[39]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[3]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[40]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[41]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[42]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[43]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[44]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[45]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[46]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[47]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[48]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[49]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[4]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[50]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[51]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[52]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[53]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[54]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[55]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[56]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[57]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[58]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[59]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[5]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[60]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[61]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[62]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[63]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[64]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[65]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[66]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[67]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[68]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[69]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[6]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[70]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[71]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[72]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[73]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[74]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[75]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[76]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[77]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[78]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[79]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[7]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[80]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[81]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[82]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[83]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[84]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[85]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[86]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[87]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[88]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[89]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[8]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[90]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[91]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[92]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[93]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[94]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[95]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[96]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[97]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[98]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[99]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[9]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[0]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[10], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[10]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[1]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[2]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[3]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[4]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[5]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[6]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[7]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[8]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[9], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[9]);
    $setuphold (posedge DRPCLK, negedge DRPDI[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[0]);
    $setuphold (posedge DRPCLK, negedge DRPDI[10], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[10]);
    $setuphold (posedge DRPCLK, negedge DRPDI[11], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[11]);
    $setuphold (posedge DRPCLK, negedge DRPDI[12], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[12]);
    $setuphold (posedge DRPCLK, negedge DRPDI[13], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[13]);
    $setuphold (posedge DRPCLK, negedge DRPDI[14], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[14]);
    $setuphold (posedge DRPCLK, negedge DRPDI[15], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[15]);
    $setuphold (posedge DRPCLK, negedge DRPDI[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[1]);
    $setuphold (posedge DRPCLK, negedge DRPDI[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[2]);
    $setuphold (posedge DRPCLK, negedge DRPDI[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[3]);
    $setuphold (posedge DRPCLK, negedge DRPDI[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[4]);
    $setuphold (posedge DRPCLK, negedge DRPDI[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[5]);
    $setuphold (posedge DRPCLK, negedge DRPDI[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[6]);
    $setuphold (posedge DRPCLK, negedge DRPDI[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[7]);
    $setuphold (posedge DRPCLK, negedge DRPDI[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[8]);
    $setuphold (posedge DRPCLK, negedge DRPDI[9], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[9]);
    $setuphold (posedge DRPCLK, negedge DRPEN, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPEN);
    $setuphold (posedge DRPCLK, negedge DRPWE, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPWE);
    $setuphold (posedge DRPCLK, posedge DRPADDR[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[0]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[10], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[10]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[1]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[2]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[3]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[4]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[5]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[6]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[7]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[8]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[9], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[9]);
    $setuphold (posedge DRPCLK, posedge DRPDI[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[0]);
    $setuphold (posedge DRPCLK, posedge DRPDI[10], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[10]);
    $setuphold (posedge DRPCLK, posedge DRPDI[11], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[11]);
    $setuphold (posedge DRPCLK, posedge DRPDI[12], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[12]);
    $setuphold (posedge DRPCLK, posedge DRPDI[13], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[13]);
    $setuphold (posedge DRPCLK, posedge DRPDI[14], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[14]);
    $setuphold (posedge DRPCLK, posedge DRPDI[15], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[15]);
    $setuphold (posedge DRPCLK, posedge DRPDI[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[1]);
    $setuphold (posedge DRPCLK, posedge DRPDI[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[2]);
    $setuphold (posedge DRPCLK, posedge DRPDI[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[3]);
    $setuphold (posedge DRPCLK, posedge DRPDI[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[4]);
    $setuphold (posedge DRPCLK, posedge DRPDI[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[5]);
    $setuphold (posedge DRPCLK, posedge DRPDI[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[6]);
    $setuphold (posedge DRPCLK, posedge DRPDI[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[7]);
    $setuphold (posedge DRPCLK, posedge DRPDI[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[8]);
    $setuphold (posedge DRPCLK, posedge DRPDI[9], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[9]);
    $setuphold (posedge DRPCLK, posedge DRPEN, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPEN);
    $setuphold (posedge DRPCLK, posedge DRPWE, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPWE);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[0]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[1]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[2]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[3]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[4]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[5]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[0]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[1]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[2]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[3]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[4]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQDONE);
    $setuphold (posedge PIPECLK, negedge PLDISABLESCRAMBLER, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDISABLESCRAMBLER);
    $setuphold (posedge PIPECLK, negedge PLEQRESETEIEOSCOUNT, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLEQRESETEIEOSCOUNT);
    $setuphold (posedge PIPECLK, negedge PLGEN3PCSDISABLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLGEN3PCSDISABLE);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[0]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[1]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[2]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[3]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[4]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[5]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[0]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[1]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[2]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[3]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[4]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQDONE);
    $setuphold (posedge PIPECLK, posedge PLDISABLESCRAMBLER, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDISABLESCRAMBLER);
    $setuphold (posedge PIPECLK, posedge PLEQRESETEIEOSCOUNT, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLEQRESETEIEOSCOUNT);
    $setuphold (posedge PIPECLK, posedge PLGEN3PCSDISABLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLGEN3PCSDISABLE);
    $setuphold (posedge RECCLK, negedge PIPERX0CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX0CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX0ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX0PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX0STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX0STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX0STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX0STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX0SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX0SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX0VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0VALID);
    $setuphold (posedge RECCLK, negedge PIPERX1CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX1CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX1ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX1PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX1STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX1STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX1STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX1STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX1SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX1SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX1VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1VALID);
    $setuphold (posedge RECCLK, negedge PIPERX2CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX2CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX2ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX2PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX2STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX2STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX2STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX2STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX2SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX2SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX2VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2VALID);
    $setuphold (posedge RECCLK, negedge PIPERX3CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX3CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX3ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX3PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX3STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX3STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX3STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX3STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX3SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX3SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX3VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3VALID);
    $setuphold (posedge RECCLK, negedge PIPERX4CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX4CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX4ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX4PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX4STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX4STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX4STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX4STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX4SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX4SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX4VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4VALID);
    $setuphold (posedge RECCLK, negedge PIPERX5CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX5CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX5ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX5PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX5STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX5STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX5STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX5STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX5SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX5SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX5VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5VALID);
    $setuphold (posedge RECCLK, negedge PIPERX6CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX6CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX6ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX6PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX6STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX6STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX6STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX6STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX6SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX6SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX6VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6VALID);
    $setuphold (posedge RECCLK, negedge PIPERX7CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX7CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX7ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX7PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX7STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX7STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX7STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX7STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX7SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX7SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX7VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7VALID);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[0]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[1]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[2]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[3]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[4]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[5]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[6]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[7]);
    $setuphold (posedge RECCLK, posedge PIPERX0CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX0CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX0ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX0PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX0STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX0STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX0STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX0STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX0SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX0SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX0VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0VALID);
    $setuphold (posedge RECCLK, posedge PIPERX1CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX1CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX1ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX1PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX1STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX1STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX1STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX1STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX1SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX1SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX1VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1VALID);
    $setuphold (posedge RECCLK, posedge PIPERX2CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX2CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX2ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX2PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX2STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX2STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX2STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX2STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX2SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX2SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX2VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2VALID);
    $setuphold (posedge RECCLK, posedge PIPERX3CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX3CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX3ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX3PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX3STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX3STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX3STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX3STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX3SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX3SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX3VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3VALID);
    $setuphold (posedge RECCLK, posedge PIPERX4CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX4CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX4ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX4PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX4STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX4STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX4STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX4STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX4SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX4SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX4VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4VALID);
    $setuphold (posedge RECCLK, posedge PIPERX5CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX5CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX5ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX5PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX5STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX5STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX5STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX5STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX5SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX5SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX5VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5VALID);
    $setuphold (posedge RECCLK, posedge PIPERX6CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX6CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX6ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX6PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX6STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX6STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX6STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX6STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX6SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX6SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX6VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6VALID);
    $setuphold (posedge RECCLK, posedge PIPERX7CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX7CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX7ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX7PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX7STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX7STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX7STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX7STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX7SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX7SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX7VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7VALID);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[0]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[1]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[2]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[3]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[4]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[5]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[6]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[7]);
    $setuphold (posedge USERCLK, negedge CFGCONFIGSPACEENABLE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGCONFIGSPACEENABLE);
    $setuphold (posedge USERCLK, negedge CFGDEVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[0]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[10]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[11]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[12]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[13]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[14]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[15]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[1]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[2]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[3]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[4]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[5]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[6]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[7]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[8]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[9]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[3]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[4]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[5]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[6]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[7]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[3]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[4]);
    $setuphold (posedge USERCLK, negedge CFGDSFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGDSFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGDSFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGDSN[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[0]);
    $setuphold (posedge USERCLK, negedge CFGDSN[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[10]);
    $setuphold (posedge USERCLK, negedge CFGDSN[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[11]);
    $setuphold (posedge USERCLK, negedge CFGDSN[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[12]);
    $setuphold (posedge USERCLK, negedge CFGDSN[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[13]);
    $setuphold (posedge USERCLK, negedge CFGDSN[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[14]);
    $setuphold (posedge USERCLK, negedge CFGDSN[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[15]);
    $setuphold (posedge USERCLK, negedge CFGDSN[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[16]);
    $setuphold (posedge USERCLK, negedge CFGDSN[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[17]);
    $setuphold (posedge USERCLK, negedge CFGDSN[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[18]);
    $setuphold (posedge USERCLK, negedge CFGDSN[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[19]);
    $setuphold (posedge USERCLK, negedge CFGDSN[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[1]);
    $setuphold (posedge USERCLK, negedge CFGDSN[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[20]);
    $setuphold (posedge USERCLK, negedge CFGDSN[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[21]);
    $setuphold (posedge USERCLK, negedge CFGDSN[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[22]);
    $setuphold (posedge USERCLK, negedge CFGDSN[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[23]);
    $setuphold (posedge USERCLK, negedge CFGDSN[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[24]);
    $setuphold (posedge USERCLK, negedge CFGDSN[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[25]);
    $setuphold (posedge USERCLK, negedge CFGDSN[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[26]);
    $setuphold (posedge USERCLK, negedge CFGDSN[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[27]);
    $setuphold (posedge USERCLK, negedge CFGDSN[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[28]);
    $setuphold (posedge USERCLK, negedge CFGDSN[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[29]);
    $setuphold (posedge USERCLK, negedge CFGDSN[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[2]);
    $setuphold (posedge USERCLK, negedge CFGDSN[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[30]);
    $setuphold (posedge USERCLK, negedge CFGDSN[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[31]);
    $setuphold (posedge USERCLK, negedge CFGDSN[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[32]);
    $setuphold (posedge USERCLK, negedge CFGDSN[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[33]);
    $setuphold (posedge USERCLK, negedge CFGDSN[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[34]);
    $setuphold (posedge USERCLK, negedge CFGDSN[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[35]);
    $setuphold (posedge USERCLK, negedge CFGDSN[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[36]);
    $setuphold (posedge USERCLK, negedge CFGDSN[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[37]);
    $setuphold (posedge USERCLK, negedge CFGDSN[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[38]);
    $setuphold (posedge USERCLK, negedge CFGDSN[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[39]);
    $setuphold (posedge USERCLK, negedge CFGDSN[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[3]);
    $setuphold (posedge USERCLK, negedge CFGDSN[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[40]);
    $setuphold (posedge USERCLK, negedge CFGDSN[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[41]);
    $setuphold (posedge USERCLK, negedge CFGDSN[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[42]);
    $setuphold (posedge USERCLK, negedge CFGDSN[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[43]);
    $setuphold (posedge USERCLK, negedge CFGDSN[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[44]);
    $setuphold (posedge USERCLK, negedge CFGDSN[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[45]);
    $setuphold (posedge USERCLK, negedge CFGDSN[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[46]);
    $setuphold (posedge USERCLK, negedge CFGDSN[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[47]);
    $setuphold (posedge USERCLK, negedge CFGDSN[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[48]);
    $setuphold (posedge USERCLK, negedge CFGDSN[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[49]);
    $setuphold (posedge USERCLK, negedge CFGDSN[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[4]);
    $setuphold (posedge USERCLK, negedge CFGDSN[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[50]);
    $setuphold (posedge USERCLK, negedge CFGDSN[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[51]);
    $setuphold (posedge USERCLK, negedge CFGDSN[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[52]);
    $setuphold (posedge USERCLK, negedge CFGDSN[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[53]);
    $setuphold (posedge USERCLK, negedge CFGDSN[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[54]);
    $setuphold (posedge USERCLK, negedge CFGDSN[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[55]);
    $setuphold (posedge USERCLK, negedge CFGDSN[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[56]);
    $setuphold (posedge USERCLK, negedge CFGDSN[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[57]);
    $setuphold (posedge USERCLK, negedge CFGDSN[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[58]);
    $setuphold (posedge USERCLK, negedge CFGDSN[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[59]);
    $setuphold (posedge USERCLK, negedge CFGDSN[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[5]);
    $setuphold (posedge USERCLK, negedge CFGDSN[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[60]);
    $setuphold (posedge USERCLK, negedge CFGDSN[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[61]);
    $setuphold (posedge USERCLK, negedge CFGDSN[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[62]);
    $setuphold (posedge USERCLK, negedge CFGDSN[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[63]);
    $setuphold (posedge USERCLK, negedge CFGDSN[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[6]);
    $setuphold (posedge USERCLK, negedge CFGDSN[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[7]);
    $setuphold (posedge USERCLK, negedge CFGDSN[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[8]);
    $setuphold (posedge USERCLK, negedge CFGDSN[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[9]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[3]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[4]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[5]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[6]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[7]);
    $setuphold (posedge USERCLK, negedge CFGERRCORIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGERRCORIN);
    $setuphold (posedge USERCLK, negedge CFGERRUNCORIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGERRUNCORIN);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATAVALID);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[0]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[10]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[11]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[12]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[13]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[14]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[15]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[16]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[17]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[18]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[19]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[1]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[20]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[21]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[22]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[23]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[24]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[25]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[26]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[27]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[28]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[29]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[2]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[30]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[31]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[3]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[4]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[5]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[6]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[7]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[8]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[9]);
    $setuphold (posedge USERCLK, negedge CFGFCSEL[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[0]);
    $setuphold (posedge USERCLK, negedge CFGFCSEL[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[1]);
    $setuphold (posedge USERCLK, negedge CFGFCSEL[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[2]);
    $setuphold (posedge USERCLK, negedge CFGFLRDONE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFLRDONE[0]);
    $setuphold (posedge USERCLK, negedge CFGFLRDONE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFLRDONE[1]);
    $setuphold (posedge USERCLK, negedge CFGHOTRESETIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGHOTRESETIN);
    $setuphold (posedge USERCLK, negedge CFGINPUTUPDATEREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINPUTUPDATEREQUEST);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIATTR[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIATTR[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIATTR[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[32]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[33]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[34]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[35]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[36]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[37]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[38]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[39]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[40]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[41]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[42]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[43]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[44]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[45]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[46]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[47]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[48]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[49]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[50]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[51]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[52]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[53]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[54]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[55]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[56]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[57]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[58]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[59]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[60]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[61]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[62]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[63]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHPRESENT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHPRESENT);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHTYPE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHTYPE[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHTYPE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHTYPE[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[32]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[33]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[34]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[35]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[36]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[37]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[38]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[39]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[40]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[41]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[42]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[43]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[44]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[45]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[46]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[47]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[48]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[49]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[50]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[51]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[52]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[53]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[54]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[55]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[56]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[57]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[58]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[59]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[60]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[61]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[62]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[63]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXINT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXINT);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTPENDING[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTPENDING[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTPENDING[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTPENDING[1]);
    $setuphold (posedge USERCLK, negedge CFGLINKTRAININGENABLE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGLINKTRAININGENABLE);
    $setuphold (posedge USERCLK, negedge CFGMCUPDATEREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMCUPDATEREQUEST);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[0]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[10]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[11]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[12]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[13]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[14]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[15]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[16]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[17]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[18]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[1]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[2]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[3]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[4]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[5]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[6]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[7]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[8]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[9]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[0]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[1]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[2]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[3]);
    $setuphold (posedge USERCLK, negedge CFGMGMTREAD, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTREAD);
    $setuphold (posedge USERCLK, negedge CFGMGMTTYPE1CFGREGACCESS, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTTYPE1CFGREGACCESS);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITE);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[0]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[10]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[11]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[12]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[13]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[14]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[15]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[16]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[17]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[18]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[19]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[1]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[20]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[21]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[22]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[23]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[24]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[25]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[26]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[27]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[28]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[29]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[2]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[30]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[31]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[3]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[4]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[5]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[6]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[7]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[8]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[9]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMIT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMIT);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[0]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[10]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[11]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[12]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[13]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[14]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[15]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[16]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[17]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[18]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[19]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[1]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[20]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[21]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[22]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[23]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[24]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[25]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[26]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[27]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[28]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[29]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[2]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[30]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[31]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[3]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[4]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[5]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[6]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[7]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[8]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[9]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITTYPE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[0]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITTYPE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[1]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITTYPE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[2]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCSTATUSCONTROL[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[0]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCSTATUSCONTROL[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[1]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCSTATUSCONTROL[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[2]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONOUTPUTREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONOUTPUTREQUEST);
    $setuphold (posedge USERCLK, negedge CFGPOWERSTATECHANGEACK, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPOWERSTATECHANGEACK);
    $setuphold (posedge USERCLK, negedge CFGREQPMTRANSITIONL23READY, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREQPMTRANSITIONL23READY);
    $setuphold (posedge USERCLK, negedge CFGREVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[0]);
    $setuphold (posedge USERCLK, negedge CFGREVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[1]);
    $setuphold (posedge USERCLK, negedge CFGREVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[2]);
    $setuphold (posedge USERCLK, negedge CFGREVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[3]);
    $setuphold (posedge USERCLK, negedge CFGREVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[4]);
    $setuphold (posedge USERCLK, negedge CFGREVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[5]);
    $setuphold (posedge USERCLK, negedge CFGREVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[6]);
    $setuphold (posedge USERCLK, negedge CFGREVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[7]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[0]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[10]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[11]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[12]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[13]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[14]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[15]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[1]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[2]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[3]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[4]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[5]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[6]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[7]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[8]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[9]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[0]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[10]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[11]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[12]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[13]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[14]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[15]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[1]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[2]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[3]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[4]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[5]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[6]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[7]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[8]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[9]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATAVALID);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[0]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[10]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[11]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[12]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[13]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[14]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[15]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[16]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[17]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[18]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[19]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[1]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[20]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[21]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[22]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[23]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[24]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[25]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[26]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[27]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[28]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[29]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[2]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[30]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[31]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[3]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[4]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[5]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[6]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[7]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[8]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[9]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[0]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[10]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[11]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[12]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[13]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[14]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[15]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[1]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[2]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[3]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[4]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[5]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[6]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[7]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[8]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[9]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[0]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[1]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[2]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[3]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[4]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[5]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[0]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[10]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[11]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[12]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[13]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[14]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[15]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[16]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[17]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[18]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[19]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[1]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[20]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[21]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[2]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[3]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[4]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[5]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[6]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[7]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[8]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[9]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[0]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[10]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[11]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[12]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[13]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[14]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[15]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[16]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[17]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[18]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[19]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[1]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[20]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[21]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[2]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[3]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[4]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[5]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[6]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[7]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[8]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[9]);
    $setuphold (posedge USERCLK, negedge PCIECQNPREQ, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_PCIECQNPREQ);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[0]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[100]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[101]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[102]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[103]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[104]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[105]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[106]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[107]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[108]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[109]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[10]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[110]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[111]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[112]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[113]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[114]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[115]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[116]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[117]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[118]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[119]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[11]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[120]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[121]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[122]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[123]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[124]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[125]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[126]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[127]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[128], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[128]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[129], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[129]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[12]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[130], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[130]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[131], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[131]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[132], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[132]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[133], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[133]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[134], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[134]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[135], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[135]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[136], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[136]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[137], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[137]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[138], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[138]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[139], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[139]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[13]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[140], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[140]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[141], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[141]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[142], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[142]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[143], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[143]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[144], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[144]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[145], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[145]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[146], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[146]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[147], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[147]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[148], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[148]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[149], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[149]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[14]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[150], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[150]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[151], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[151]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[152], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[152]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[153], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[153]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[154], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[154]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[155], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[155]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[156], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[156]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[157], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[157]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[158], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[158]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[159], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[159]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[15]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[160], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[160]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[161], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[161]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[162], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[162]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[163], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[163]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[164], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[164]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[165], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[165]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[166], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[166]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[167], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[167]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[168], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[168]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[169], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[169]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[16]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[170], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[170]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[171], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[171]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[172], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[172]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[173], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[173]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[174], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[174]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[175], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[175]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[176], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[176]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[177], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[177]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[178], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[178]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[179], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[179]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[17]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[180], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[180]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[181], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[181]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[182], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[182]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[183], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[183]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[184], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[184]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[185], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[185]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[186], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[186]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[187], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[187]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[188], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[188]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[189], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[189]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[18]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[190], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[190]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[191], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[191]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[192], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[192]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[193], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[193]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[194], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[194]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[195], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[195]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[196], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[196]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[197], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[197]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[198], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[198]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[199], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[199]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[19]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[1]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[200], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[200]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[201], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[201]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[202], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[202]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[203], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[203]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[204], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[204]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[205], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[205]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[206], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[206]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[207], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[207]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[208], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[208]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[209], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[209]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[20]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[210], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[210]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[211], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[211]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[212], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[212]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[213], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[213]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[214], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[214]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[215], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[215]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[216], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[216]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[217], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[217]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[218], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[218]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[219], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[219]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[21]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[220], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[220]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[221], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[221]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[222], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[222]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[223], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[223]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[224], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[224]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[225], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[225]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[226], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[226]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[227], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[227]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[228], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[228]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[229], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[229]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[22]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[230], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[230]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[231], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[231]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[232], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[232]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[233], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[233]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[234], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[234]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[235], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[235]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[236], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[236]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[237], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[237]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[238], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[238]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[239], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[239]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[23]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[240], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[240]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[241], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[241]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[242], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[242]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[243], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[243]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[244], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[244]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[245], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[245]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[246], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[246]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[247], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[247]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[248], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[248]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[249], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[249]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[24]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[250], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[250]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[251], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[251]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[252], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[252]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[253], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[253]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[254], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[254]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[255], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[255]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[25]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[26]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[27]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[28]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[29]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[2]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[30]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[31]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[32]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[33]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[34]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[35]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[36]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[37]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[38]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[39]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[3]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[40]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[41]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[42]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[43]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[44]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[45]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[46]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[47]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[48]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[49]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[4]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[50]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[51]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[52]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[53]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[54]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[55]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[56]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[57]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[58]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[59]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[5]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[60]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[61]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[62]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[63]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[64]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[65]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[66]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[67]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[68]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[69]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[6]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[70]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[71]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[72]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[73]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[74]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[75]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[76]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[77]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[78]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[79]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[7]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[80]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[81]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[82]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[83]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[84]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[85]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[86]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[87]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[88]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[89]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[8]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[90]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[91]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[92]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[93]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[94]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[95]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[96]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[97]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[98]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[99]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[9]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[0]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[1]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[2]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[3]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[4]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[5]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[6]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[7]);
    $setuphold (posedge USERCLK, negedge SAXISCCTLAST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTLAST);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[0]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[10]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[11]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[12]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[13]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[14]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[15]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[16]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[17]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[18]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[19]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[1]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[20]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[21]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[22]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[23]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[24]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[25]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[26]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[27]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[28]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[29]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[2]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[30]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[31]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[32]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[3]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[4]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[5]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[6]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[7]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[8]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[9]);
    $setuphold (posedge USERCLK, negedge SAXISCCTVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTVALID);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[0]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[100]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[101]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[102]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[103]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[104]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[105]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[106]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[107]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[108]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[109]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[10]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[110]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[111]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[112]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[113]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[114]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[115]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[116]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[117]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[118]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[119]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[11]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[120]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[121]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[122]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[123]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[124]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[125]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[126]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[127]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[128], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[128]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[129], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[129]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[12]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[130], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[130]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[131], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[131]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[132], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[132]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[133], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[133]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[134], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[134]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[135], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[135]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[136], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[136]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[137], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[137]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[138], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[138]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[139], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[139]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[13]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[140], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[140]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[141], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[141]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[142], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[142]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[143], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[143]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[144], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[144]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[145], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[145]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[146], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[146]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[147], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[147]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[148], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[148]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[149], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[149]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[14]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[150], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[150]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[151], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[151]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[152], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[152]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[153], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[153]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[154], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[154]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[155], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[155]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[156], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[156]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[157], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[157]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[158], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[158]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[159], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[159]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[15]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[160], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[160]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[161], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[161]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[162], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[162]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[163], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[163]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[164], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[164]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[165], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[165]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[166], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[166]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[167], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[167]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[168], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[168]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[169], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[169]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[16]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[170], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[170]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[171], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[171]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[172], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[172]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[173], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[173]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[174], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[174]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[175], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[175]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[176], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[176]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[177], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[177]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[178], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[178]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[179], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[179]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[17]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[180], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[180]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[181], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[181]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[182], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[182]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[183], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[183]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[184], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[184]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[185], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[185]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[186], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[186]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[187], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[187]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[188], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[188]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[189], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[189]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[18]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[190], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[190]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[191], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[191]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[192], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[192]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[193], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[193]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[194], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[194]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[195], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[195]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[196], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[196]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[197], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[197]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[198], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[198]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[199], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[199]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[19]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[1]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[200], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[200]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[201], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[201]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[202], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[202]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[203], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[203]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[204], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[204]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[205], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[205]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[206], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[206]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[207], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[207]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[208], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[208]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[209], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[209]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[20]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[210], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[210]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[211], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[211]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[212], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[212]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[213], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[213]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[214], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[214]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[215], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[215]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[216], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[216]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[217], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[217]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[218], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[218]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[219], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[219]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[21]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[220], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[220]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[221], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[221]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[222], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[222]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[223], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[223]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[224], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[224]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[225], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[225]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[226], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[226]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[227], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[227]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[228], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[228]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[229], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[229]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[22]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[230], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[230]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[231], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[231]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[232], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[232]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[233], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[233]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[234], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[234]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[235], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[235]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[236], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[236]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[237], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[237]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[238], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[238]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[239], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[239]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[23]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[240], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[240]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[241], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[241]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[242], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[242]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[243], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[243]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[244], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[244]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[245], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[245]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[246], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[246]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[247], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[247]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[248], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[248]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[249], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[249]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[24]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[250], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[250]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[251], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[251]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[252], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[252]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[253], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[253]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[254], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[254]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[255], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[255]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[25]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[26]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[27]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[28]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[29]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[2]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[30]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[31]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[32]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[33]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[34]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[35]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[36]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[37]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[38]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[39]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[3]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[40]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[41]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[42]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[43]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[44]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[45]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[46]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[47]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[48]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[49]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[4]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[50]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[51]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[52]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[53]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[54]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[55]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[56]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[57]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[58]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[59]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[5]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[60]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[61]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[62]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[63]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[64]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[65]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[66]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[67]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[68]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[69]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[6]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[70]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[71]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[72]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[73]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[74]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[75]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[76]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[77]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[78]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[79]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[7]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[80]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[81]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[82]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[83]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[84]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[85]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[86]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[87]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[88]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[89]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[8]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[90]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[91]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[92]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[93]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[94]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[95]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[96]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[97]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[98]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[99]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[9]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[0]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[1]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[2]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[3]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[4]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[5]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[6]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[7]);
    $setuphold (posedge USERCLK, negedge SAXISRQTLAST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTLAST);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[0]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[10]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[11]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[12]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[13]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[14]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[15]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[16]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[17]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[18]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[19]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[1]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[20]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[21]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[22]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[23]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[24]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[25]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[26]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[27]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[28]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[29]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[2]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[30]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[31]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[32]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[33]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[34]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[35]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[36]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[37]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[38]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[39]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[3]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[40]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[41]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[42]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[43]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[44]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[45]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[46]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[47]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[48]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[49]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[4]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[50]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[51]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[52]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[53]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[54]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[55]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[56]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[57]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[58]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[59]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[5]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[6]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[7]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[8]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[9]);
    $setuphold (posedge USERCLK, negedge SAXISRQTVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTVALID);
    $setuphold (posedge USERCLK, posedge CFGCONFIGSPACEENABLE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGCONFIGSPACEENABLE);
    $setuphold (posedge USERCLK, posedge CFGDEVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[0]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[10]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[11]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[12]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[13]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[14]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[15]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[1]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[2]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[3]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[4]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[5]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[6]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[7]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[8]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[9]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[3]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[4]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[5]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[6]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[7]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[3]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[4]);
    $setuphold (posedge USERCLK, posedge CFGDSFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGDSFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGDSFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGDSN[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[0]);
    $setuphold (posedge USERCLK, posedge CFGDSN[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[10]);
    $setuphold (posedge USERCLK, posedge CFGDSN[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[11]);
    $setuphold (posedge USERCLK, posedge CFGDSN[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[12]);
    $setuphold (posedge USERCLK, posedge CFGDSN[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[13]);
    $setuphold (posedge USERCLK, posedge CFGDSN[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[14]);
    $setuphold (posedge USERCLK, posedge CFGDSN[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[15]);
    $setuphold (posedge USERCLK, posedge CFGDSN[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[16]);
    $setuphold (posedge USERCLK, posedge CFGDSN[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[17]);
    $setuphold (posedge USERCLK, posedge CFGDSN[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[18]);
    $setuphold (posedge USERCLK, posedge CFGDSN[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[19]);
    $setuphold (posedge USERCLK, posedge CFGDSN[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[1]);
    $setuphold (posedge USERCLK, posedge CFGDSN[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[20]);
    $setuphold (posedge USERCLK, posedge CFGDSN[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[21]);
    $setuphold (posedge USERCLK, posedge CFGDSN[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[22]);
    $setuphold (posedge USERCLK, posedge CFGDSN[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[23]);
    $setuphold (posedge USERCLK, posedge CFGDSN[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[24]);
    $setuphold (posedge USERCLK, posedge CFGDSN[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[25]);
    $setuphold (posedge USERCLK, posedge CFGDSN[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[26]);
    $setuphold (posedge USERCLK, posedge CFGDSN[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[27]);
    $setuphold (posedge USERCLK, posedge CFGDSN[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[28]);
    $setuphold (posedge USERCLK, posedge CFGDSN[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[29]);
    $setuphold (posedge USERCLK, posedge CFGDSN[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[2]);
    $setuphold (posedge USERCLK, posedge CFGDSN[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[30]);
    $setuphold (posedge USERCLK, posedge CFGDSN[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[31]);
    $setuphold (posedge USERCLK, posedge CFGDSN[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[32]);
    $setuphold (posedge USERCLK, posedge CFGDSN[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[33]);
    $setuphold (posedge USERCLK, posedge CFGDSN[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[34]);
    $setuphold (posedge USERCLK, posedge CFGDSN[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[35]);
    $setuphold (posedge USERCLK, posedge CFGDSN[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[36]);
    $setuphold (posedge USERCLK, posedge CFGDSN[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[37]);
    $setuphold (posedge USERCLK, posedge CFGDSN[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[38]);
    $setuphold (posedge USERCLK, posedge CFGDSN[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[39]);
    $setuphold (posedge USERCLK, posedge CFGDSN[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[3]);
    $setuphold (posedge USERCLK, posedge CFGDSN[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[40]);
    $setuphold (posedge USERCLK, posedge CFGDSN[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[41]);
    $setuphold (posedge USERCLK, posedge CFGDSN[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[42]);
    $setuphold (posedge USERCLK, posedge CFGDSN[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[43]);
    $setuphold (posedge USERCLK, posedge CFGDSN[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[44]);
    $setuphold (posedge USERCLK, posedge CFGDSN[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[45]);
    $setuphold (posedge USERCLK, posedge CFGDSN[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[46]);
    $setuphold (posedge USERCLK, posedge CFGDSN[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[47]);
    $setuphold (posedge USERCLK, posedge CFGDSN[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[48]);
    $setuphold (posedge USERCLK, posedge CFGDSN[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[49]);
    $setuphold (posedge USERCLK, posedge CFGDSN[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[4]);
    $setuphold (posedge USERCLK, posedge CFGDSN[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[50]);
    $setuphold (posedge USERCLK, posedge CFGDSN[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[51]);
    $setuphold (posedge USERCLK, posedge CFGDSN[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[52]);
    $setuphold (posedge USERCLK, posedge CFGDSN[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[53]);
    $setuphold (posedge USERCLK, posedge CFGDSN[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[54]);
    $setuphold (posedge USERCLK, posedge CFGDSN[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[55]);
    $setuphold (posedge USERCLK, posedge CFGDSN[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[56]);
    $setuphold (posedge USERCLK, posedge CFGDSN[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[57]);
    $setuphold (posedge USERCLK, posedge CFGDSN[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[58]);
    $setuphold (posedge USERCLK, posedge CFGDSN[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[59]);
    $setuphold (posedge USERCLK, posedge CFGDSN[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[5]);
    $setuphold (posedge USERCLK, posedge CFGDSN[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[60]);
    $setuphold (posedge USERCLK, posedge CFGDSN[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[61]);
    $setuphold (posedge USERCLK, posedge CFGDSN[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[62]);
    $setuphold (posedge USERCLK, posedge CFGDSN[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[63]);
    $setuphold (posedge USERCLK, posedge CFGDSN[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[6]);
    $setuphold (posedge USERCLK, posedge CFGDSN[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[7]);
    $setuphold (posedge USERCLK, posedge CFGDSN[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[8]);
    $setuphold (posedge USERCLK, posedge CFGDSN[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[9]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[3]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[4]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[5]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[6]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[7]);
    $setuphold (posedge USERCLK, posedge CFGERRCORIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGERRCORIN);
    $setuphold (posedge USERCLK, posedge CFGERRUNCORIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGERRUNCORIN);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATAVALID);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[0]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[10]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[11]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[12]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[13]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[14]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[15]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[16]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[17]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[18]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[19]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[1]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[20]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[21]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[22]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[23]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[24]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[25]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[26]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[27]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[28]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[29]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[2]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[30]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[31]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[3]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[4]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[5]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[6]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[7]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[8]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[9]);
    $setuphold (posedge USERCLK, posedge CFGFCSEL[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[0]);
    $setuphold (posedge USERCLK, posedge CFGFCSEL[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[1]);
    $setuphold (posedge USERCLK, posedge CFGFCSEL[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[2]);
    $setuphold (posedge USERCLK, posedge CFGFLRDONE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFLRDONE[0]);
    $setuphold (posedge USERCLK, posedge CFGFLRDONE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFLRDONE[1]);
    $setuphold (posedge USERCLK, posedge CFGHOTRESETIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGHOTRESETIN);
    $setuphold (posedge USERCLK, posedge CFGINPUTUPDATEREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINPUTUPDATEREQUEST);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIATTR[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIATTR[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIATTR[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[32]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[33]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[34]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[35]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[36]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[37]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[38]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[39]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[40]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[41]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[42]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[43]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[44]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[45]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[46]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[47]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[48]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[49]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[50]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[51]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[52]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[53]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[54]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[55]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[56]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[57]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[58]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[59]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[60]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[61]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[62]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[63]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHPRESENT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHPRESENT);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHTYPE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHTYPE[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHTYPE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHTYPE[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[32]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[33]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[34]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[35]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[36]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[37]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[38]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[39]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[40]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[41]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[42]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[43]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[44]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[45]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[46]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[47]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[48]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[49]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[50]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[51]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[52]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[53]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[54]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[55]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[56]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[57]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[58]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[59]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[60]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[61]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[62]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[63]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXINT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXINT);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTPENDING[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTPENDING[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTPENDING[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTPENDING[1]);
    $setuphold (posedge USERCLK, posedge CFGLINKTRAININGENABLE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGLINKTRAININGENABLE);
    $setuphold (posedge USERCLK, posedge CFGMCUPDATEREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMCUPDATEREQUEST);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[0]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[10]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[11]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[12]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[13]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[14]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[15]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[16]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[17]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[18]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[1]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[2]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[3]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[4]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[5]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[6]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[7]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[8]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[9]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[0]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[1]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[2]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[3]);
    $setuphold (posedge USERCLK, posedge CFGMGMTREAD, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTREAD);
    $setuphold (posedge USERCLK, posedge CFGMGMTTYPE1CFGREGACCESS, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTTYPE1CFGREGACCESS);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITE);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[0]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[10]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[11]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[12]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[13]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[14]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[15]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[16]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[17]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[18]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[19]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[1]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[20]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[21]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[22]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[23]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[24]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[25]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[26]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[27]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[28]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[29]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[2]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[30]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[31]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[3]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[4]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[5]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[6]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[7]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[8]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[9]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMIT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMIT);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[0]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[10]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[11]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[12]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[13]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[14]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[15]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[16]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[17]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[18]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[19]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[1]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[20]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[21]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[22]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[23]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[24]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[25]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[26]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[27]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[28]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[29]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[2]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[30]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[31]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[3]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[4]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[5]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[6]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[7]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[8]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[9]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITTYPE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[0]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITTYPE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[1]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITTYPE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[2]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCSTATUSCONTROL[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[0]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCSTATUSCONTROL[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[1]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCSTATUSCONTROL[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[2]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONOUTPUTREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONOUTPUTREQUEST);
    $setuphold (posedge USERCLK, posedge CFGPOWERSTATECHANGEACK, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPOWERSTATECHANGEACK);
    $setuphold (posedge USERCLK, posedge CFGREQPMTRANSITIONL23READY, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREQPMTRANSITIONL23READY);
    $setuphold (posedge USERCLK, posedge CFGREVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[0]);
    $setuphold (posedge USERCLK, posedge CFGREVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[1]);
    $setuphold (posedge USERCLK, posedge CFGREVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[2]);
    $setuphold (posedge USERCLK, posedge CFGREVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[3]);
    $setuphold (posedge USERCLK, posedge CFGREVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[4]);
    $setuphold (posedge USERCLK, posedge CFGREVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[5]);
    $setuphold (posedge USERCLK, posedge CFGREVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[6]);
    $setuphold (posedge USERCLK, posedge CFGREVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[7]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[0]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[10]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[11]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[12]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[13]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[14]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[15]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[1]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[2]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[3]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[4]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[5]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[6]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[7]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[8]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[9]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[0]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[10]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[11]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[12]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[13]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[14]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[15]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[1]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[2]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[3]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[4]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[5]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[6]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[7]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[8]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[9]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATAVALID);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[0]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[10]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[11]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[12]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[13]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[14]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[15]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[16]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[17]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[18]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[19]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[1]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[20]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[21]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[22]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[23]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[24]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[25]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[26]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[27]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[28]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[29]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[2]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[30]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[31]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[3]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[4]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[5]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[6]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[7]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[8]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[9]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[0]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[10]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[11]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[12]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[13]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[14]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[15]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[1]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[2]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[3]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[4]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[5]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[6]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[7]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[8]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[9]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[0]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[1]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[2]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[3]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[4]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[5]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[0]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[10]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[11]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[12]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[13]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[14]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[15]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[16]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[17]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[18]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[19]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[1]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[20]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[21]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[2]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[3]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[4]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[5]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[6]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[7]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[8]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[9]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[0]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[10]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[11]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[12]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[13]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[14]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[15]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[16]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[17]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[18]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[19]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[1]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[20]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[21]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[2]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[3]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[4]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[5]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[6]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[7]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[8]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[9]);
    $setuphold (posedge USERCLK, posedge PCIECQNPREQ, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_PCIECQNPREQ);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[0]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[100]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[101]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[102]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[103]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[104]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[105]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[106]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[107]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[108]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[109]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[10]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[110]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[111]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[112]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[113]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[114]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[115]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[116]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[117]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[118]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[119]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[11]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[120]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[121]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[122]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[123]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[124]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[125]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[126]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[127]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[128], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[128]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[129], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[129]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[12]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[130], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[130]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[131], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[131]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[132], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[132]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[133], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[133]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[134], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[134]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[135], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[135]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[136], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[136]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[137], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[137]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[138], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[138]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[139], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[139]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[13]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[140], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[140]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[141], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[141]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[142], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[142]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[143], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[143]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[144], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[144]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[145], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[145]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[146], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[146]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[147], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[147]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[148], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[148]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[149], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[149]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[14]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[150], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[150]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[151], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[151]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[152], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[152]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[153], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[153]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[154], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[154]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[155], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[155]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[156], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[156]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[157], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[157]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[158], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[158]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[159], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[159]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[15]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[160], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[160]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[161], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[161]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[162], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[162]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[163], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[163]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[164], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[164]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[165], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[165]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[166], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[166]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[167], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[167]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[168], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[168]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[169], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[169]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[16]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[170], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[170]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[171], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[171]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[172], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[172]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[173], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[173]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[174], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[174]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[175], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[175]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[176], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[176]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[177], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[177]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[178], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[178]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[179], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[179]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[17]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[180], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[180]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[181], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[181]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[182], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[182]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[183], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[183]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[184], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[184]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[185], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[185]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[186], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[186]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[187], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[187]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[188], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[188]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[189], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[189]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[18]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[190], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[190]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[191], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[191]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[192], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[192]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[193], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[193]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[194], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[194]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[195], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[195]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[196], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[196]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[197], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[197]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[198], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[198]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[199], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[199]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[19]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[1]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[200], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[200]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[201], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[201]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[202], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[202]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[203], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[203]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[204], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[204]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[205], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[205]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[206], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[206]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[207], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[207]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[208], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[208]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[209], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[209]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[20]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[210], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[210]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[211], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[211]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[212], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[212]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[213], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[213]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[214], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[214]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[215], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[215]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[216], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[216]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[217], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[217]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[218], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[218]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[219], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[219]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[21]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[220], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[220]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[221], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[221]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[222], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[222]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[223], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[223]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[224], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[224]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[225], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[225]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[226], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[226]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[227], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[227]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[228], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[228]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[229], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[229]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[22]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[230], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[230]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[231], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[231]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[232], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[232]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[233], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[233]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[234], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[234]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[235], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[235]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[236], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[236]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[237], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[237]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[238], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[238]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[239], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[239]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[23]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[240], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[240]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[241], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[241]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[242], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[242]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[243], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[243]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[244], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[244]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[245], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[245]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[246], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[246]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[247], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[247]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[248], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[248]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[249], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[249]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[24]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[250], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[250]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[251], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[251]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[252], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[252]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[253], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[253]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[254], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[254]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[255], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[255]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[25]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[26]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[27]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[28]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[29]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[2]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[30]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[31]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[32]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[33]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[34]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[35]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[36]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[37]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[38]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[39]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[3]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[40]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[41]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[42]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[43]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[44]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[45]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[46]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[47]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[48]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[49]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[4]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[50]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[51]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[52]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[53]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[54]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[55]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[56]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[57]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[58]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[59]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[5]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[60]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[61]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[62]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[63]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[64]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[65]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[66]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[67]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[68]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[69]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[6]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[70]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[71]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[72]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[73]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[74]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[75]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[76]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[77]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[78]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[79]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[7]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[80]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[81]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[82]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[83]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[84]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[85]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[86]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[87]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[88]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[89]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[8]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[90]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[91]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[92]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[93]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[94]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[95]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[96]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[97]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[98]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[99]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[9]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[0]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[1]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[2]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[3]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[4]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[5]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[6]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[7]);
    $setuphold (posedge USERCLK, posedge SAXISCCTLAST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTLAST);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[0]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[10]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[11]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[12]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[13]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[14]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[15]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[16]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[17]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[18]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[19]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[1]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[20]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[21]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[22]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[23]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[24]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[25]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[26]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[27]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[28]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[29]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[2]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[30]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[31]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[32]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[3]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[4]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[5]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[6]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[7]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[8]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[9]);
    $setuphold (posedge USERCLK, posedge SAXISCCTVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTVALID);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[0]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[100]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[101]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[102]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[103]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[104]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[105]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[106]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[107]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[108]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[109]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[10]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[110]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[111]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[112]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[113]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[114]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[115]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[116]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[117]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[118]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[119]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[11]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[120]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[121]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[122]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[123]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[124]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[125]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[126]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[127]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[128], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[128]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[129], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[129]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[12]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[130], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[130]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[131], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[131]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[132], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[132]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[133], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[133]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[134], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[134]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[135], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[135]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[136], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[136]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[137], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[137]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[138], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[138]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[139], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[139]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[13]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[140], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[140]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[141], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[141]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[142], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[142]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[143], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[143]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[144], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[144]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[145], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[145]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[146], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[146]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[147], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[147]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[148], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[148]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[149], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[149]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[14]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[150], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[150]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[151], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[151]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[152], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[152]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[153], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[153]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[154], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[154]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[155], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[155]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[156], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[156]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[157], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[157]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[158], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[158]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[159], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[159]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[15]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[160], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[160]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[161], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[161]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[162], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[162]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[163], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[163]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[164], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[164]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[165], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[165]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[166], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[166]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[167], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[167]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[168], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[168]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[169], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[169]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[16]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[170], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[170]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[171], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[171]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[172], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[172]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[173], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[173]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[174], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[174]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[175], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[175]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[176], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[176]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[177], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[177]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[178], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[178]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[179], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[179]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[17]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[180], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[180]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[181], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[181]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[182], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[182]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[183], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[183]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[184], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[184]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[185], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[185]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[186], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[186]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[187], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[187]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[188], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[188]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[189], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[189]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[18]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[190], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[190]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[191], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[191]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[192], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[192]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[193], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[193]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[194], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[194]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[195], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[195]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[196], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[196]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[197], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[197]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[198], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[198]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[199], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[199]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[19]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[1]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[200], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[200]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[201], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[201]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[202], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[202]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[203], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[203]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[204], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[204]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[205], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[205]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[206], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[206]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[207], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[207]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[208], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[208]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[209], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[209]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[20]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[210], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[210]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[211], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[211]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[212], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[212]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[213], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[213]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[214], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[214]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[215], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[215]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[216], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[216]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[217], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[217]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[218], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[218]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[219], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[219]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[21]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[220], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[220]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[221], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[221]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[222], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[222]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[223], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[223]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[224], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[224]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[225], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[225]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[226], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[226]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[227], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[227]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[228], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[228]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[229], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[229]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[22]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[230], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[230]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[231], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[231]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[232], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[232]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[233], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[233]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[234], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[234]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[235], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[235]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[236], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[236]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[237], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[237]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[238], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[238]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[239], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[239]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[23]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[240], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[240]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[241], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[241]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[242], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[242]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[243], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[243]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[244], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[244]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[245], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[245]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[246], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[246]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[247], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[247]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[248], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[248]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[249], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[249]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[24]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[250], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[250]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[251], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[251]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[252], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[252]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[253], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[253]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[254], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[254]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[255], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[255]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[25]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[26]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[27]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[28]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[29]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[2]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[30]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[31]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[32]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[33]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[34]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[35]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[36]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[37]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[38]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[39]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[3]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[40]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[41]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[42]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[43]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[44]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[45]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[46]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[47]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[48]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[49]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[4]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[50]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[51]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[52]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[53]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[54]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[55]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[56]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[57]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[58]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[59]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[5]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[60]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[61]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[62]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[63]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[64]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[65]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[66]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[67]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[68]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[69]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[6]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[70]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[71]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[72]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[73]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[74]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[75]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[76]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[77]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[78]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[79]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[7]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[80]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[81]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[82]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[83]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[84]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[85]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[86]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[87]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[88]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[89]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[8]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[90]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[91]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[92]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[93]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[94]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[95]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[96]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[97]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[98]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[99]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[9]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[0]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[1]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[2]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[3]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[4]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[5]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[6]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[7]);
    $setuphold (posedge USERCLK, posedge SAXISRQTLAST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTLAST);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[0]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[10]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[11]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[12]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[13]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[14]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[15]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[16]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[17]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[18]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[19]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[1]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[20]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[21]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[22]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[23]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[24]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[25]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[26]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[27]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[28]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[29]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[2]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[30]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[31]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[32]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[33]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[34]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[35]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[36]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[37]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[38]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[39]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[3]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[40]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[41]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[42]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[43]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[44]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[45]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[46]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[47]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[48]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[49]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[4]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[50]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[51]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[52]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[53]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[54]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[55]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[56]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[57]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[58]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[59]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[5]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[6]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[7]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[8]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[9]);
    $setuphold (posedge USERCLK, posedge SAXISRQTVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTVALID);
`endif

    ( CORECLK *> DBGDATAOUT[0]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[10]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[11]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[12]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[13]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[14]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[15]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[1]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[2]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[3]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[4]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[5]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[6]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[7]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[8]) = (0, 0);
    ( CORECLK *> DBGDATAOUT[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[4]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[5]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[6]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[7]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[8]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[4]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[5]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[6]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[7]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[8]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADENABLEL[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADENABLEL[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADENABLEL[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADENABLEL[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[4]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[5]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[6]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[7]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[8]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[4]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[5]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[6]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[7]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[8]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[10]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[11]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[12]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[13]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[14]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[15]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[16]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[17]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[18]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[19]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[20]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[21]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[22]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[23]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[24]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[25]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[26]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[27]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[28]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[29]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[30]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[31]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[32]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[33]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[34]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[35]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[36]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[37]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[38]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[39]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[40]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[41]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[42]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[43]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[44]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[45]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[46]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[47]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[48]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[49]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[4]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[50]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[51]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[52]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[53]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[54]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[55]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[56]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[57]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[58]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[59]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[5]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[60]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[61]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[62]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[63]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[64]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[65]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[66]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[67]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[68]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[69]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[6]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[70]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[71]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[7]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[8]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEENABLEL[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEENABLEL[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEENABLEL[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEENABLEL[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[4]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[5]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[6]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[7]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[8]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[4]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[5]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[6]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[7]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[8]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADENABLEU[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADENABLEU[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADENABLEU[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADENABLEU[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[4]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[5]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[6]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[7]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[8]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[4]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[5]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[6]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[7]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[8]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[10]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[11]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[12]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[13]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[14]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[15]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[16]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[17]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[18]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[19]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[20]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[21]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[22]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[23]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[24]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[25]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[26]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[27]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[28]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[29]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[30]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[31]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[32]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[33]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[34]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[35]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[36]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[37]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[38]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[39]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[3]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[40]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[41]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[42]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[43]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[44]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[45]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[46]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[47]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[48]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[49]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[4]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[50]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[51]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[52]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[53]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[54]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[55]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[56]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[57]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[58]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[59]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[5]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[60]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[61]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[62]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[63]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[64]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[65]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[66]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[67]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[68]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[69]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[6]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[70]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[71]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[7]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[8]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[9]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEENABLEU[0]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEENABLEU[1]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEENABLEU[2]) = (0, 0);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEENABLEU[3]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[0]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[1]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[2]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[3]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[4]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[5]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[6]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[7]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[8]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMREADENABLE[0]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMREADENABLE[1]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[0]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[100]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[101]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[102]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[103]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[104]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[105]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[106]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[107]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[108]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[109]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[10]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[110]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[111]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[112]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[113]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[114]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[115]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[116]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[117]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[118]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[119]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[11]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[120]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[121]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[122]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[123]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[124]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[125]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[126]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[127]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[128]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[129]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[12]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[130]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[131]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[132]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[133]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[134]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[135]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[136]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[137]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[138]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[139]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[13]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[140]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[141]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[142]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[143]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[14]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[15]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[16]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[17]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[18]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[19]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[1]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[20]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[21]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[22]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[23]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[24]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[25]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[26]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[27]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[28]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[29]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[2]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[30]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[31]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[32]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[33]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[34]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[35]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[36]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[37]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[38]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[39]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[3]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[40]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[41]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[42]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[43]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[44]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[45]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[46]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[47]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[48]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[49]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[4]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[50]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[51]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[52]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[53]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[54]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[55]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[56]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[57]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[58]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[59]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[5]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[60]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[61]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[62]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[63]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[64]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[65]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[66]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[67]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[68]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[69]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[6]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[70]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[71]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[72]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[73]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[74]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[75]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[76]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[77]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[78]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[79]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[7]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[80]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[81]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[82]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[83]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[84]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[85]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[86]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[87]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[88]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[89]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[8]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[90]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[91]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[92]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[93]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[94]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[95]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[96]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[97]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[98]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[99]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[9]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEENABLE[0]) = (0, 0);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEENABLE[1]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[0]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[1]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[2]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[3]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[4]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[5]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[6]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[7]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[8]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[0]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[1]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[2]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[3]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[4]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[5]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[6]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[7]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[8]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADENABLE[0]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADENABLE[1]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADENABLE[2]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADENABLE[3]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[0]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[1]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[2]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[3]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[4]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[5]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[6]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[7]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[8]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[0]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[1]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[2]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[3]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[4]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[5]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[6]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[7]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[8]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[0]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[100]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[101]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[102]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[103]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[104]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[105]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[106]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[107]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[108]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[109]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[10]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[110]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[111]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[112]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[113]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[114]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[115]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[116]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[117]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[118]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[119]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[11]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[120]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[121]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[122]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[123]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[124]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[125]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[126]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[127]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[128]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[129]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[12]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[130]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[131]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[132]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[133]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[134]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[135]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[136]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[137]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[138]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[139]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[13]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[140]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[141]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[142]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[143]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[14]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[15]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[16]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[17]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[18]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[19]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[1]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[20]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[21]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[22]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[23]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[24]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[25]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[26]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[27]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[28]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[29]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[2]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[30]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[31]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[32]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[33]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[34]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[35]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[36]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[37]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[38]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[39]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[3]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[40]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[41]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[42]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[43]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[44]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[45]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[46]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[47]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[48]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[49]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[4]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[50]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[51]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[52]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[53]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[54]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[55]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[56]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[57]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[58]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[59]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[5]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[60]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[61]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[62]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[63]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[64]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[65]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[66]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[67]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[68]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[69]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[6]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[70]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[71]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[72]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[73]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[74]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[75]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[76]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[77]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[78]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[79]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[7]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[80]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[81]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[82]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[83]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[84]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[85]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[86]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[87]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[88]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[89]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[8]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[90]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[91]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[92]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[93]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[94]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[95]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[96]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[97]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[98]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[99]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[9]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEENABLE[0]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEENABLE[1]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEENABLE[2]) = (0, 0);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEENABLE[3]) = (0, 0);
    ( DRPCLK *> DRPDO[0]) = (0, 0);
    ( DRPCLK *> DRPDO[10]) = (0, 0);
    ( DRPCLK *> DRPDO[11]) = (0, 0);
    ( DRPCLK *> DRPDO[12]) = (0, 0);
    ( DRPCLK *> DRPDO[13]) = (0, 0);
    ( DRPCLK *> DRPDO[14]) = (0, 0);
    ( DRPCLK *> DRPDO[15]) = (0, 0);
    ( DRPCLK *> DRPDO[1]) = (0, 0);
    ( DRPCLK *> DRPDO[2]) = (0, 0);
    ( DRPCLK *> DRPDO[3]) = (0, 0);
    ( DRPCLK *> DRPDO[4]) = (0, 0);
    ( DRPCLK *> DRPDO[5]) = (0, 0);
    ( DRPCLK *> DRPDO[6]) = (0, 0);
    ( DRPCLK *> DRPDO[7]) = (0, 0);
    ( DRPCLK *> DRPDO[8]) = (0, 0);
    ( DRPCLK *> DRPDO[9]) = (0, 0);
    ( DRPCLK *> DRPRDY) = (0, 0);
    ( PIPECLK *> PIPERX0EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPERX0EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPERX0EQLPLFFS[0]) = (0, 0);
    ( PIPECLK *> PIPERX0EQLPLFFS[1]) = (0, 0);
    ( PIPECLK *> PIPERX0EQLPLFFS[2]) = (0, 0);
    ( PIPECLK *> PIPERX0EQLPLFFS[3]) = (0, 0);
    ( PIPECLK *> PIPERX0EQLPLFFS[4]) = (0, 0);
    ( PIPECLK *> PIPERX0EQLPLFFS[5]) = (0, 0);
    ( PIPECLK *> PIPERX0EQLPTXPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX0EQLPTXPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX0EQLPTXPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX0EQLPTXPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPERX0EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX0EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX0EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX0POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX1EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPERX1EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPERX1EQLPLFFS[0]) = (0, 0);
    ( PIPECLK *> PIPERX1EQLPLFFS[1]) = (0, 0);
    ( PIPECLK *> PIPERX1EQLPLFFS[2]) = (0, 0);
    ( PIPECLK *> PIPERX1EQLPLFFS[3]) = (0, 0);
    ( PIPECLK *> PIPERX1EQLPLFFS[4]) = (0, 0);
    ( PIPECLK *> PIPERX1EQLPLFFS[5]) = (0, 0);
    ( PIPECLK *> PIPERX1EQLPTXPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX1EQLPTXPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX1EQLPTXPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX1EQLPTXPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPERX1EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX1EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX1EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX1POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX2EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPERX2EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPERX2EQLPLFFS[0]) = (0, 0);
    ( PIPECLK *> PIPERX2EQLPLFFS[1]) = (0, 0);
    ( PIPECLK *> PIPERX2EQLPLFFS[2]) = (0, 0);
    ( PIPECLK *> PIPERX2EQLPLFFS[3]) = (0, 0);
    ( PIPECLK *> PIPERX2EQLPLFFS[4]) = (0, 0);
    ( PIPECLK *> PIPERX2EQLPLFFS[5]) = (0, 0);
    ( PIPECLK *> PIPERX2EQLPTXPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX2EQLPTXPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX2EQLPTXPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX2EQLPTXPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPERX2EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX2EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX2EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX2POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX3EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPERX3EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPERX3EQLPLFFS[0]) = (0, 0);
    ( PIPECLK *> PIPERX3EQLPLFFS[1]) = (0, 0);
    ( PIPECLK *> PIPERX3EQLPLFFS[2]) = (0, 0);
    ( PIPECLK *> PIPERX3EQLPLFFS[3]) = (0, 0);
    ( PIPECLK *> PIPERX3EQLPLFFS[4]) = (0, 0);
    ( PIPECLK *> PIPERX3EQLPLFFS[5]) = (0, 0);
    ( PIPECLK *> PIPERX3EQLPTXPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX3EQLPTXPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX3EQLPTXPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX3EQLPTXPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPERX3EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX3EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX3EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX3POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX4EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPERX4EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPERX4EQLPLFFS[0]) = (0, 0);
    ( PIPECLK *> PIPERX4EQLPLFFS[1]) = (0, 0);
    ( PIPECLK *> PIPERX4EQLPLFFS[2]) = (0, 0);
    ( PIPECLK *> PIPERX4EQLPLFFS[3]) = (0, 0);
    ( PIPECLK *> PIPERX4EQLPLFFS[4]) = (0, 0);
    ( PIPECLK *> PIPERX4EQLPLFFS[5]) = (0, 0);
    ( PIPECLK *> PIPERX4EQLPTXPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX4EQLPTXPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX4EQLPTXPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX4EQLPTXPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPERX4EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX4EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX4EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX4POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX5EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPERX5EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPERX5EQLPLFFS[0]) = (0, 0);
    ( PIPECLK *> PIPERX5EQLPLFFS[1]) = (0, 0);
    ( PIPECLK *> PIPERX5EQLPLFFS[2]) = (0, 0);
    ( PIPECLK *> PIPERX5EQLPLFFS[3]) = (0, 0);
    ( PIPECLK *> PIPERX5EQLPLFFS[4]) = (0, 0);
    ( PIPECLK *> PIPERX5EQLPLFFS[5]) = (0, 0);
    ( PIPECLK *> PIPERX5EQLPTXPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX5EQLPTXPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX5EQLPTXPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX5EQLPTXPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPERX5EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX5EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX5EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX5POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX6EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPERX6EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPERX6EQLPLFFS[0]) = (0, 0);
    ( PIPECLK *> PIPERX6EQLPLFFS[1]) = (0, 0);
    ( PIPECLK *> PIPERX6EQLPLFFS[2]) = (0, 0);
    ( PIPECLK *> PIPERX6EQLPLFFS[3]) = (0, 0);
    ( PIPECLK *> PIPERX6EQLPLFFS[4]) = (0, 0);
    ( PIPECLK *> PIPERX6EQLPLFFS[5]) = (0, 0);
    ( PIPECLK *> PIPERX6EQLPTXPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX6EQLPTXPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX6EQLPTXPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX6EQLPTXPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPERX6EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX6EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX6EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX6POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX7EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPERX7EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPERX7EQLPLFFS[0]) = (0, 0);
    ( PIPECLK *> PIPERX7EQLPLFFS[1]) = (0, 0);
    ( PIPECLK *> PIPERX7EQLPLFFS[2]) = (0, 0);
    ( PIPECLK *> PIPERX7EQLPLFFS[3]) = (0, 0);
    ( PIPECLK *> PIPERX7EQLPLFFS[4]) = (0, 0);
    ( PIPECLK *> PIPERX7EQLPLFFS[5]) = (0, 0);
    ( PIPECLK *> PIPERX7EQLPTXPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX7EQLPTXPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX7EQLPTXPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX7EQLPTXPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPERX7EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPERX7EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPERX7EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPERX7POLARITY) = (0, 0);
    ( PIPECLK *> PIPETX0CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX0CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX0COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX0DATAVALID) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[16]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[17]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[18]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[19]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[20]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[21]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[22]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[23]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[24]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[25]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[26]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[27]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[28]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[29]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[30]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[31]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX0ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX0EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPETX0EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPETX0EQDEEMPH[0]) = (0, 0);
    ( PIPECLK *> PIPETX0EQDEEMPH[1]) = (0, 0);
    ( PIPECLK *> PIPETX0EQDEEMPH[2]) = (0, 0);
    ( PIPECLK *> PIPETX0EQDEEMPH[3]) = (0, 0);
    ( PIPECLK *> PIPETX0EQDEEMPH[4]) = (0, 0);
    ( PIPECLK *> PIPETX0EQDEEMPH[5]) = (0, 0);
    ( PIPECLK *> PIPETX0EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPETX0EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPETX0EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPETX0EQPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPETX0POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX0POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX0STARTBLOCK) = (0, 0);
    ( PIPECLK *> PIPETX0SYNCHEADER[0]) = (0, 0);
    ( PIPECLK *> PIPETX0SYNCHEADER[1]) = (0, 0);
    ( PIPECLK *> PIPETX1CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX1CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX1COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX1DATAVALID) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[16]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[17]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[18]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[19]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[20]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[21]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[22]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[23]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[24]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[25]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[26]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[27]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[28]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[29]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[30]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[31]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX1ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX1EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPETX1EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPETX1EQDEEMPH[0]) = (0, 0);
    ( PIPECLK *> PIPETX1EQDEEMPH[1]) = (0, 0);
    ( PIPECLK *> PIPETX1EQDEEMPH[2]) = (0, 0);
    ( PIPECLK *> PIPETX1EQDEEMPH[3]) = (0, 0);
    ( PIPECLK *> PIPETX1EQDEEMPH[4]) = (0, 0);
    ( PIPECLK *> PIPETX1EQDEEMPH[5]) = (0, 0);
    ( PIPECLK *> PIPETX1EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPETX1EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPETX1EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPETX1EQPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPETX1POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX1POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX1STARTBLOCK) = (0, 0);
    ( PIPECLK *> PIPETX1SYNCHEADER[0]) = (0, 0);
    ( PIPECLK *> PIPETX1SYNCHEADER[1]) = (0, 0);
    ( PIPECLK *> PIPETX2CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX2CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX2COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX2DATAVALID) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[16]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[17]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[18]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[19]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[20]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[21]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[22]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[23]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[24]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[25]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[26]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[27]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[28]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[29]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[30]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[31]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX2ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX2EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPETX2EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPETX2EQDEEMPH[0]) = (0, 0);
    ( PIPECLK *> PIPETX2EQDEEMPH[1]) = (0, 0);
    ( PIPECLK *> PIPETX2EQDEEMPH[2]) = (0, 0);
    ( PIPECLK *> PIPETX2EQDEEMPH[3]) = (0, 0);
    ( PIPECLK *> PIPETX2EQDEEMPH[4]) = (0, 0);
    ( PIPECLK *> PIPETX2EQDEEMPH[5]) = (0, 0);
    ( PIPECLK *> PIPETX2EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPETX2EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPETX2EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPETX2EQPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPETX2POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX2POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX2STARTBLOCK) = (0, 0);
    ( PIPECLK *> PIPETX2SYNCHEADER[0]) = (0, 0);
    ( PIPECLK *> PIPETX2SYNCHEADER[1]) = (0, 0);
    ( PIPECLK *> PIPETX3CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX3CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX3COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX3DATAVALID) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[16]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[17]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[18]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[19]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[20]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[21]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[22]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[23]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[24]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[25]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[26]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[27]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[28]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[29]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[30]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[31]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX3ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX3EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPETX3EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPETX3EQDEEMPH[0]) = (0, 0);
    ( PIPECLK *> PIPETX3EQDEEMPH[1]) = (0, 0);
    ( PIPECLK *> PIPETX3EQDEEMPH[2]) = (0, 0);
    ( PIPECLK *> PIPETX3EQDEEMPH[3]) = (0, 0);
    ( PIPECLK *> PIPETX3EQDEEMPH[4]) = (0, 0);
    ( PIPECLK *> PIPETX3EQDEEMPH[5]) = (0, 0);
    ( PIPECLK *> PIPETX3EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPETX3EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPETX3EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPETX3EQPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPETX3POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX3POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX3STARTBLOCK) = (0, 0);
    ( PIPECLK *> PIPETX3SYNCHEADER[0]) = (0, 0);
    ( PIPECLK *> PIPETX3SYNCHEADER[1]) = (0, 0);
    ( PIPECLK *> PIPETX4CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX4CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX4COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX4DATAVALID) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[16]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[17]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[18]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[19]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[20]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[21]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[22]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[23]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[24]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[25]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[26]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[27]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[28]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[29]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[30]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[31]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX4ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX4EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPETX4EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPETX4EQDEEMPH[0]) = (0, 0);
    ( PIPECLK *> PIPETX4EQDEEMPH[1]) = (0, 0);
    ( PIPECLK *> PIPETX4EQDEEMPH[2]) = (0, 0);
    ( PIPECLK *> PIPETX4EQDEEMPH[3]) = (0, 0);
    ( PIPECLK *> PIPETX4EQDEEMPH[4]) = (0, 0);
    ( PIPECLK *> PIPETX4EQDEEMPH[5]) = (0, 0);
    ( PIPECLK *> PIPETX4EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPETX4EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPETX4EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPETX4EQPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPETX4POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX4POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX4STARTBLOCK) = (0, 0);
    ( PIPECLK *> PIPETX4SYNCHEADER[0]) = (0, 0);
    ( PIPECLK *> PIPETX4SYNCHEADER[1]) = (0, 0);
    ( PIPECLK *> PIPETX5CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX5CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX5COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX5DATAVALID) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[16]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[17]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[18]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[19]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[20]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[21]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[22]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[23]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[24]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[25]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[26]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[27]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[28]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[29]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[30]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[31]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX5ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX5EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPETX5EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPETX5EQDEEMPH[0]) = (0, 0);
    ( PIPECLK *> PIPETX5EQDEEMPH[1]) = (0, 0);
    ( PIPECLK *> PIPETX5EQDEEMPH[2]) = (0, 0);
    ( PIPECLK *> PIPETX5EQDEEMPH[3]) = (0, 0);
    ( PIPECLK *> PIPETX5EQDEEMPH[4]) = (0, 0);
    ( PIPECLK *> PIPETX5EQDEEMPH[5]) = (0, 0);
    ( PIPECLK *> PIPETX5EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPETX5EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPETX5EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPETX5EQPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPETX5POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX5POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX5STARTBLOCK) = (0, 0);
    ( PIPECLK *> PIPETX5SYNCHEADER[0]) = (0, 0);
    ( PIPECLK *> PIPETX5SYNCHEADER[1]) = (0, 0);
    ( PIPECLK *> PIPETX6CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX6CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX6COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX6DATAVALID) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[16]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[17]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[18]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[19]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[20]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[21]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[22]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[23]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[24]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[25]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[26]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[27]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[28]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[29]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[30]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[31]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX6ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX6EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPETX6EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPETX6EQDEEMPH[0]) = (0, 0);
    ( PIPECLK *> PIPETX6EQDEEMPH[1]) = (0, 0);
    ( PIPECLK *> PIPETX6EQDEEMPH[2]) = (0, 0);
    ( PIPECLK *> PIPETX6EQDEEMPH[3]) = (0, 0);
    ( PIPECLK *> PIPETX6EQDEEMPH[4]) = (0, 0);
    ( PIPECLK *> PIPETX6EQDEEMPH[5]) = (0, 0);
    ( PIPECLK *> PIPETX6EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPETX6EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPETX6EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPETX6EQPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPETX6POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX6POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX6STARTBLOCK) = (0, 0);
    ( PIPECLK *> PIPETX6SYNCHEADER[0]) = (0, 0);
    ( PIPECLK *> PIPETX6SYNCHEADER[1]) = (0, 0);
    ( PIPECLK *> PIPETX7CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX7CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX7COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX7DATAVALID) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[16]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[17]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[18]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[19]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[20]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[21]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[22]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[23]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[24]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[25]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[26]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[27]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[28]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[29]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[30]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[31]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX7ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX7EQCONTROL[0]) = (0, 0);
    ( PIPECLK *> PIPETX7EQCONTROL[1]) = (0, 0);
    ( PIPECLK *> PIPETX7EQDEEMPH[0]) = (0, 0);
    ( PIPECLK *> PIPETX7EQDEEMPH[1]) = (0, 0);
    ( PIPECLK *> PIPETX7EQDEEMPH[2]) = (0, 0);
    ( PIPECLK *> PIPETX7EQDEEMPH[3]) = (0, 0);
    ( PIPECLK *> PIPETX7EQDEEMPH[4]) = (0, 0);
    ( PIPECLK *> PIPETX7EQDEEMPH[5]) = (0, 0);
    ( PIPECLK *> PIPETX7EQPRESET[0]) = (0, 0);
    ( PIPECLK *> PIPETX7EQPRESET[1]) = (0, 0);
    ( PIPECLK *> PIPETX7EQPRESET[2]) = (0, 0);
    ( PIPECLK *> PIPETX7EQPRESET[3]) = (0, 0);
    ( PIPECLK *> PIPETX7POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX7POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX7STARTBLOCK) = (0, 0);
    ( PIPECLK *> PIPETX7SYNCHEADER[0]) = (0, 0);
    ( PIPECLK *> PIPETX7SYNCHEADER[1]) = (0, 0);
    ( PIPECLK *> PIPETXDEEMPH) = (0, 0);
    ( PIPECLK *> PIPETXMARGIN[0]) = (0, 0);
    ( PIPECLK *> PIPETXMARGIN[1]) = (0, 0);
    ( PIPECLK *> PIPETXMARGIN[2]) = (0, 0);
    ( PIPECLK *> PIPETXRATE[0]) = (0, 0);
    ( PIPECLK *> PIPETXRATE[1]) = (0, 0);
    ( PIPECLK *> PIPETXRCVRDET) = (0, 0);
    ( PIPECLK *> PIPETXRESET) = (0, 0);
    ( PIPECLK *> PIPETXSWING) = (0, 0);
    ( PIPECLK *> PLEQINPROGRESS) = (0, 0);
    ( PIPECLK *> PLEQPHASE[0]) = (0, 0);
    ( PIPECLK *> PLEQPHASE[1]) = (0, 0);
    ( RECCLK *> PLGEN3PCSRXSLIDE[0]) = (0, 0);
    ( RECCLK *> PLGEN3PCSRXSLIDE[1]) = (0, 0);
    ( RECCLK *> PLGEN3PCSRXSLIDE[2]) = (0, 0);
    ( RECCLK *> PLGEN3PCSRXSLIDE[3]) = (0, 0);
    ( RECCLK *> PLGEN3PCSRXSLIDE[4]) = (0, 0);
    ( RECCLK *> PLGEN3PCSRXSLIDE[5]) = (0, 0);
    ( RECCLK *> PLGEN3PCSRXSLIDE[6]) = (0, 0);
    ( RECCLK *> PLGEN3PCSRXSLIDE[7]) = (0, 0);
    ( USERCLK *> CFGCURRENTSPEED[0]) = (0, 0);
    ( USERCLK *> CFGCURRENTSPEED[1]) = (0, 0);
    ( USERCLK *> CFGCURRENTSPEED[2]) = (0, 0);
    ( USERCLK *> CFGDPASUBSTATECHANGE[0]) = (0, 0);
    ( USERCLK *> CFGDPASUBSTATECHANGE[1]) = (0, 0);
    ( USERCLK *> CFGERRCOROUT) = (0, 0);
    ( USERCLK *> CFGERRFATALOUT) = (0, 0);
    ( USERCLK *> CFGERRNONFATALOUT) = (0, 0);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[0]) = (0, 0);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[1]) = (0, 0);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[2]) = (0, 0);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[3]) = (0, 0);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[4]) = (0, 0);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[5]) = (0, 0);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[6]) = (0, 0);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[7]) = (0, 0);
    ( USERCLK *> CFGEXTREADRECEIVED) = (0, 0);
    ( USERCLK *> CFGEXTREGISTERNUMBER[0]) = (0, 0);
    ( USERCLK *> CFGEXTREGISTERNUMBER[1]) = (0, 0);
    ( USERCLK *> CFGEXTREGISTERNUMBER[2]) = (0, 0);
    ( USERCLK *> CFGEXTREGISTERNUMBER[3]) = (0, 0);
    ( USERCLK *> CFGEXTREGISTERNUMBER[4]) = (0, 0);
    ( USERCLK *> CFGEXTREGISTERNUMBER[5]) = (0, 0);
    ( USERCLK *> CFGEXTREGISTERNUMBER[6]) = (0, 0);
    ( USERCLK *> CFGEXTREGISTERNUMBER[7]) = (0, 0);
    ( USERCLK *> CFGEXTREGISTERNUMBER[8]) = (0, 0);
    ( USERCLK *> CFGEXTREGISTERNUMBER[9]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEBYTEENABLE[0]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEBYTEENABLE[1]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEBYTEENABLE[2]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEBYTEENABLE[3]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[0]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[10]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[11]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[12]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[13]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[14]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[15]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[16]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[17]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[18]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[19]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[1]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[20]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[21]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[22]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[23]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[24]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[25]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[26]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[27]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[28]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[29]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[2]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[30]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[31]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[3]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[4]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[5]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[6]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[7]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[8]) = (0, 0);
    ( USERCLK *> CFGEXTWRITEDATA[9]) = (0, 0);
    ( USERCLK *> CFGEXTWRITERECEIVED) = (0, 0);
    ( USERCLK *> CFGFCCPLD[0]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[10]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[11]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[1]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[2]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[3]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[4]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[5]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[6]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[7]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[8]) = (0, 0);
    ( USERCLK *> CFGFCCPLD[9]) = (0, 0);
    ( USERCLK *> CFGFCCPLH[0]) = (0, 0);
    ( USERCLK *> CFGFCCPLH[1]) = (0, 0);
    ( USERCLK *> CFGFCCPLH[2]) = (0, 0);
    ( USERCLK *> CFGFCCPLH[3]) = (0, 0);
    ( USERCLK *> CFGFCCPLH[4]) = (0, 0);
    ( USERCLK *> CFGFCCPLH[5]) = (0, 0);
    ( USERCLK *> CFGFCCPLH[6]) = (0, 0);
    ( USERCLK *> CFGFCCPLH[7]) = (0, 0);
    ( USERCLK *> CFGFCNPD[0]) = (0, 0);
    ( USERCLK *> CFGFCNPD[10]) = (0, 0);
    ( USERCLK *> CFGFCNPD[11]) = (0, 0);
    ( USERCLK *> CFGFCNPD[1]) = (0, 0);
    ( USERCLK *> CFGFCNPD[2]) = (0, 0);
    ( USERCLK *> CFGFCNPD[3]) = (0, 0);
    ( USERCLK *> CFGFCNPD[4]) = (0, 0);
    ( USERCLK *> CFGFCNPD[5]) = (0, 0);
    ( USERCLK *> CFGFCNPD[6]) = (0, 0);
    ( USERCLK *> CFGFCNPD[7]) = (0, 0);
    ( USERCLK *> CFGFCNPD[8]) = (0, 0);
    ( USERCLK *> CFGFCNPD[9]) = (0, 0);
    ( USERCLK *> CFGFCNPH[0]) = (0, 0);
    ( USERCLK *> CFGFCNPH[1]) = (0, 0);
    ( USERCLK *> CFGFCNPH[2]) = (0, 0);
    ( USERCLK *> CFGFCNPH[3]) = (0, 0);
    ( USERCLK *> CFGFCNPH[4]) = (0, 0);
    ( USERCLK *> CFGFCNPH[5]) = (0, 0);
    ( USERCLK *> CFGFCNPH[6]) = (0, 0);
    ( USERCLK *> CFGFCNPH[7]) = (0, 0);
    ( USERCLK *> CFGFCPD[0]) = (0, 0);
    ( USERCLK *> CFGFCPD[10]) = (0, 0);
    ( USERCLK *> CFGFCPD[11]) = (0, 0);
    ( USERCLK *> CFGFCPD[1]) = (0, 0);
    ( USERCLK *> CFGFCPD[2]) = (0, 0);
    ( USERCLK *> CFGFCPD[3]) = (0, 0);
    ( USERCLK *> CFGFCPD[4]) = (0, 0);
    ( USERCLK *> CFGFCPD[5]) = (0, 0);
    ( USERCLK *> CFGFCPD[6]) = (0, 0);
    ( USERCLK *> CFGFCPD[7]) = (0, 0);
    ( USERCLK *> CFGFCPD[8]) = (0, 0);
    ( USERCLK *> CFGFCPD[9]) = (0, 0);
    ( USERCLK *> CFGFCPH[0]) = (0, 0);
    ( USERCLK *> CFGFCPH[1]) = (0, 0);
    ( USERCLK *> CFGFCPH[2]) = (0, 0);
    ( USERCLK *> CFGFCPH[3]) = (0, 0);
    ( USERCLK *> CFGFCPH[4]) = (0, 0);
    ( USERCLK *> CFGFCPH[5]) = (0, 0);
    ( USERCLK *> CFGFCPH[6]) = (0, 0);
    ( USERCLK *> CFGFCPH[7]) = (0, 0);
    ( USERCLK *> CFGFLRINPROCESS[0]) = (0, 0);
    ( USERCLK *> CFGFLRINPROCESS[1]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[0]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[1]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[2]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[3]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[4]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[5]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONSTATUS[0]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONSTATUS[1]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONSTATUS[2]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONSTATUS[3]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONSTATUS[4]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONSTATUS[5]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONSTATUS[6]) = (0, 0);
    ( USERCLK *> CFGFUNCTIONSTATUS[7]) = (0, 0);
    ( USERCLK *> CFGHOTRESETOUT) = (0, 0);
    ( USERCLK *> CFGINPUTUPDATEDONE) = (0, 0);
    ( USERCLK *> CFGINTERRUPTAOUTPUT) = (0, 0);
    ( USERCLK *> CFGINTERRUPTBOUTPUT) = (0, 0);
    ( USERCLK *> CFGINTERRUPTCOUTPUT) = (0, 0);
    ( USERCLK *> CFGINTERRUPTDOUTPUT) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[0]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[10]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[11]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[12]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[13]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[14]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[15]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[16]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[17]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[18]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[19]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[1]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[20]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[21]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[22]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[23]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[24]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[25]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[26]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[27]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[28]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[29]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[2]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[30]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[31]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[3]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[4]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[5]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[6]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[7]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[8]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIDATA[9]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIENABLE[0]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIENABLE[1]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIFAIL) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIMASKUPDATE) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[0]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[1]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[2]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[3]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[4]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[5]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSISENT) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[0]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[1]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[2]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[3]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[4]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[5]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXENABLE[0]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXENABLE[1]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXFAIL) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXMASK[0]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXMASK[1]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXSENT) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[0]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[1]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[2]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[3]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[4]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[5]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[0]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[1]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[2]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[3]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[4]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[5]) = (0, 0);
    ( USERCLK *> CFGINTERRUPTSENT) = (0, 0);
    ( USERCLK *> CFGLINKPOWERSTATE[0]) = (0, 0);
    ( USERCLK *> CFGLINKPOWERSTATE[1]) = (0, 0);
    ( USERCLK *> CFGLOCALERROR) = (0, 0);
    ( USERCLK *> CFGLTRENABLE) = (0, 0);
    ( USERCLK *> CFGLTSSMSTATE[0]) = (0, 0);
    ( USERCLK *> CFGLTSSMSTATE[1]) = (0, 0);
    ( USERCLK *> CFGLTSSMSTATE[2]) = (0, 0);
    ( USERCLK *> CFGLTSSMSTATE[3]) = (0, 0);
    ( USERCLK *> CFGLTSSMSTATE[4]) = (0, 0);
    ( USERCLK *> CFGLTSSMSTATE[5]) = (0, 0);
    ( USERCLK *> CFGMAXPAYLOAD[0]) = (0, 0);
    ( USERCLK *> CFGMAXPAYLOAD[1]) = (0, 0);
    ( USERCLK *> CFGMAXPAYLOAD[2]) = (0, 0);
    ( USERCLK *> CFGMAXREADREQ[0]) = (0, 0);
    ( USERCLK *> CFGMAXREADREQ[1]) = (0, 0);
    ( USERCLK *> CFGMAXREADREQ[2]) = (0, 0);
    ( USERCLK *> CFGMCUPDATEDONE) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[0]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[10]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[11]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[12]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[13]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[14]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[15]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[16]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[17]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[18]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[19]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[1]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[20]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[21]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[22]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[23]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[24]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[25]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[26]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[27]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[28]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[29]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[2]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[30]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[31]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[3]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[4]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[5]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[6]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[7]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[8]) = (0, 0);
    ( USERCLK *> CFGMGMTREADDATA[9]) = (0, 0);
    ( USERCLK *> CFGMGMTREADWRITEDONE) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVED) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDDATA[0]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDDATA[1]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDDATA[2]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDDATA[3]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDDATA[4]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDDATA[5]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDDATA[6]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDDATA[7]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDTYPE[0]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDTYPE[1]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDTYPE[2]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDTYPE[3]) = (0, 0);
    ( USERCLK *> CFGMSGRECEIVEDTYPE[4]) = (0, 0);
    ( USERCLK *> CFGMSGTRANSMITDONE) = (0, 0);
    ( USERCLK *> CFGNEGOTIATEDWIDTH[0]) = (0, 0);
    ( USERCLK *> CFGNEGOTIATEDWIDTH[1]) = (0, 0);
    ( USERCLK *> CFGNEGOTIATEDWIDTH[2]) = (0, 0);
    ( USERCLK *> CFGNEGOTIATEDWIDTH[3]) = (0, 0);
    ( USERCLK *> CFGOBFFENABLE[0]) = (0, 0);
    ( USERCLK *> CFGOBFFENABLE[1]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[0]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[10]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[11]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[12]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[13]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[14]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[15]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[1]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[2]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[3]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[4]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[5]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[6]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[7]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[8]) = (0, 0);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[9]) = (0, 0);
    ( USERCLK *> CFGPERFUNCTIONUPDATEDONE) = (0, 0);
    ( USERCLK *> CFGPHYLINKDOWN) = (0, 0);
    ( USERCLK *> CFGPHYLINKSTATUS[0]) = (0, 0);
    ( USERCLK *> CFGPHYLINKSTATUS[1]) = (0, 0);
    ( USERCLK *> CFGPLSTATUSCHANGE) = (0, 0);
    ( USERCLK *> CFGPOWERSTATECHANGEINTERRUPT) = (0, 0);
    ( USERCLK *> CFGRCBSTATUS[0]) = (0, 0);
    ( USERCLK *> CFGRCBSTATUS[1]) = (0, 0);
    ( USERCLK *> CFGTPHFUNCTIONNUM[0]) = (0, 0);
    ( USERCLK *> CFGTPHFUNCTIONNUM[1]) = (0, 0);
    ( USERCLK *> CFGTPHFUNCTIONNUM[2]) = (0, 0);
    ( USERCLK *> CFGTPHREQUESTERENABLE[0]) = (0, 0);
    ( USERCLK *> CFGTPHREQUESTERENABLE[1]) = (0, 0);
    ( USERCLK *> CFGTPHSTMODE[0]) = (0, 0);
    ( USERCLK *> CFGTPHSTMODE[1]) = (0, 0);
    ( USERCLK *> CFGTPHSTMODE[2]) = (0, 0);
    ( USERCLK *> CFGTPHSTMODE[3]) = (0, 0);
    ( USERCLK *> CFGTPHSTMODE[4]) = (0, 0);
    ( USERCLK *> CFGTPHSTMODE[5]) = (0, 0);
    ( USERCLK *> CFGTPHSTTADDRESS[0]) = (0, 0);
    ( USERCLK *> CFGTPHSTTADDRESS[1]) = (0, 0);
    ( USERCLK *> CFGTPHSTTADDRESS[2]) = (0, 0);
    ( USERCLK *> CFGTPHSTTADDRESS[3]) = (0, 0);
    ( USERCLK *> CFGTPHSTTADDRESS[4]) = (0, 0);
    ( USERCLK *> CFGTPHSTTREADENABLE) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEBYTEVALID[0]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEBYTEVALID[1]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEBYTEVALID[2]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEBYTEVALID[3]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[0]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[10]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[11]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[12]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[13]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[14]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[15]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[16]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[17]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[18]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[19]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[1]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[20]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[21]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[22]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[23]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[24]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[25]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[26]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[27]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[28]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[29]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[2]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[30]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[31]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[3]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[4]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[5]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[6]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[7]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[8]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEDATA[9]) = (0, 0);
    ( USERCLK *> CFGTPHSTTWRITEENABLE) = (0, 0);
    ( USERCLK *> CFGVFFLRINPROCESS[0]) = (0, 0);
    ( USERCLK *> CFGVFFLRINPROCESS[1]) = (0, 0);
    ( USERCLK *> CFGVFFLRINPROCESS[2]) = (0, 0);
    ( USERCLK *> CFGVFFLRINPROCESS[3]) = (0, 0);
    ( USERCLK *> CFGVFFLRINPROCESS[4]) = (0, 0);
    ( USERCLK *> CFGVFFLRINPROCESS[5]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[0]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[10]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[11]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[12]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[13]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[14]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[15]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[16]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[17]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[1]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[2]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[3]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[4]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[5]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[6]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[7]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[8]) = (0, 0);
    ( USERCLK *> CFGVFPOWERSTATE[9]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[0]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[10]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[11]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[1]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[2]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[3]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[4]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[5]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[6]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[7]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[8]) = (0, 0);
    ( USERCLK *> CFGVFSTATUS[9]) = (0, 0);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[0]) = (0, 0);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[1]) = (0, 0);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[2]) = (0, 0);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[3]) = (0, 0);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[4]) = (0, 0);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[5]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[0]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[10]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[11]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[12]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[13]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[14]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[15]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[16]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[17]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[1]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[2]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[3]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[4]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[5]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[6]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[7]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[8]) = (0, 0);
    ( USERCLK *> CFGVFTPHSTMODE[9]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[0]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[100]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[101]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[102]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[103]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[104]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[105]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[106]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[107]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[108]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[109]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[10]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[110]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[111]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[112]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[113]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[114]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[115]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[116]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[117]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[118]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[119]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[11]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[120]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[121]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[122]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[123]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[124]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[125]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[126]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[127]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[128]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[129]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[12]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[130]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[131]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[132]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[133]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[134]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[135]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[136]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[137]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[138]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[139]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[13]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[140]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[141]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[142]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[143]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[144]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[145]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[146]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[147]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[148]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[149]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[14]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[150]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[151]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[152]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[153]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[154]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[155]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[156]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[157]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[158]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[159]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[15]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[160]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[161]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[162]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[163]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[164]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[165]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[166]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[167]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[168]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[169]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[16]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[170]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[171]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[172]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[173]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[174]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[175]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[176]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[177]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[178]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[179]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[17]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[180]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[181]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[182]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[183]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[184]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[185]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[186]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[187]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[188]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[189]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[18]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[190]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[191]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[192]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[193]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[194]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[195]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[196]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[197]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[198]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[199]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[19]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[1]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[200]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[201]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[202]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[203]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[204]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[205]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[206]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[207]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[208]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[209]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[20]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[210]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[211]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[212]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[213]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[214]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[215]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[216]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[217]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[218]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[219]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[21]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[220]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[221]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[222]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[223]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[224]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[225]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[226]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[227]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[228]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[229]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[22]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[230]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[231]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[232]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[233]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[234]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[235]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[236]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[237]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[238]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[239]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[23]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[240]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[241]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[242]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[243]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[244]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[245]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[246]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[247]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[248]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[249]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[24]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[250]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[251]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[252]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[253]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[254]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[255]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[25]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[26]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[27]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[28]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[29]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[2]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[30]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[31]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[32]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[33]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[34]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[35]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[36]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[37]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[38]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[39]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[3]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[40]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[41]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[42]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[43]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[44]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[45]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[46]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[47]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[48]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[49]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[4]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[50]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[51]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[52]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[53]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[54]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[55]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[56]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[57]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[58]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[59]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[5]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[60]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[61]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[62]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[63]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[64]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[65]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[66]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[67]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[68]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[69]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[6]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[70]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[71]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[72]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[73]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[74]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[75]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[76]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[77]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[78]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[79]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[7]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[80]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[81]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[82]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[83]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[84]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[85]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[86]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[87]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[88]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[89]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[8]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[90]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[91]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[92]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[93]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[94]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[95]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[96]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[97]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[98]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[99]) = (0, 0);
    ( USERCLK *> MAXISCQTDATA[9]) = (0, 0);
    ( USERCLK *> MAXISCQTKEEP[0]) = (0, 0);
    ( USERCLK *> MAXISCQTKEEP[1]) = (0, 0);
    ( USERCLK *> MAXISCQTKEEP[2]) = (0, 0);
    ( USERCLK *> MAXISCQTKEEP[3]) = (0, 0);
    ( USERCLK *> MAXISCQTKEEP[4]) = (0, 0);
    ( USERCLK *> MAXISCQTKEEP[5]) = (0, 0);
    ( USERCLK *> MAXISCQTKEEP[6]) = (0, 0);
    ( USERCLK *> MAXISCQTKEEP[7]) = (0, 0);
    ( USERCLK *> MAXISCQTLAST) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[0]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[10]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[11]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[12]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[13]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[14]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[15]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[16]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[17]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[18]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[19]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[1]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[20]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[21]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[22]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[23]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[24]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[25]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[26]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[27]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[28]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[29]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[2]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[30]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[31]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[32]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[33]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[34]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[35]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[36]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[37]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[38]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[39]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[3]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[40]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[41]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[42]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[43]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[44]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[45]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[46]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[47]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[48]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[49]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[4]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[50]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[51]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[52]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[53]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[54]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[55]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[56]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[57]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[58]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[59]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[5]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[60]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[61]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[62]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[63]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[64]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[65]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[66]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[67]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[68]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[69]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[6]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[70]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[71]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[72]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[73]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[74]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[75]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[76]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[77]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[78]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[79]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[7]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[80]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[81]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[82]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[83]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[84]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[8]) = (0, 0);
    ( USERCLK *> MAXISCQTUSER[9]) = (0, 0);
    ( USERCLK *> MAXISCQTVALID) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[0]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[100]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[101]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[102]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[103]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[104]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[105]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[106]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[107]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[108]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[109]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[10]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[110]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[111]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[112]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[113]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[114]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[115]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[116]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[117]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[118]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[119]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[11]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[120]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[121]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[122]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[123]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[124]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[125]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[126]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[127]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[128]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[129]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[12]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[130]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[131]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[132]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[133]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[134]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[135]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[136]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[137]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[138]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[139]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[13]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[140]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[141]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[142]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[143]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[144]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[145]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[146]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[147]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[148]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[149]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[14]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[150]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[151]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[152]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[153]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[154]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[155]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[156]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[157]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[158]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[159]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[15]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[160]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[161]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[162]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[163]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[164]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[165]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[166]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[167]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[168]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[169]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[16]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[170]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[171]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[172]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[173]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[174]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[175]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[176]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[177]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[178]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[179]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[17]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[180]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[181]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[182]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[183]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[184]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[185]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[186]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[187]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[188]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[189]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[18]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[190]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[191]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[192]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[193]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[194]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[195]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[196]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[197]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[198]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[199]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[19]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[1]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[200]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[201]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[202]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[203]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[204]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[205]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[206]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[207]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[208]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[209]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[20]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[210]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[211]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[212]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[213]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[214]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[215]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[216]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[217]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[218]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[219]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[21]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[220]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[221]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[222]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[223]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[224]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[225]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[226]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[227]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[228]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[229]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[22]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[230]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[231]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[232]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[233]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[234]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[235]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[236]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[237]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[238]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[239]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[23]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[240]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[241]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[242]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[243]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[244]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[245]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[246]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[247]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[248]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[249]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[24]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[250]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[251]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[252]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[253]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[254]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[255]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[25]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[26]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[27]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[28]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[29]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[2]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[30]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[31]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[32]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[33]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[34]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[35]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[36]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[37]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[38]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[39]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[3]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[40]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[41]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[42]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[43]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[44]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[45]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[46]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[47]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[48]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[49]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[4]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[50]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[51]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[52]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[53]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[54]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[55]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[56]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[57]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[58]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[59]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[5]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[60]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[61]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[62]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[63]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[64]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[65]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[66]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[67]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[68]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[69]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[6]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[70]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[71]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[72]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[73]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[74]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[75]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[76]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[77]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[78]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[79]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[7]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[80]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[81]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[82]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[83]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[84]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[85]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[86]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[87]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[88]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[89]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[8]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[90]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[91]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[92]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[93]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[94]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[95]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[96]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[97]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[98]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[99]) = (0, 0);
    ( USERCLK *> MAXISRCTDATA[9]) = (0, 0);
    ( USERCLK *> MAXISRCTKEEP[0]) = (0, 0);
    ( USERCLK *> MAXISRCTKEEP[1]) = (0, 0);
    ( USERCLK *> MAXISRCTKEEP[2]) = (0, 0);
    ( USERCLK *> MAXISRCTKEEP[3]) = (0, 0);
    ( USERCLK *> MAXISRCTKEEP[4]) = (0, 0);
    ( USERCLK *> MAXISRCTKEEP[5]) = (0, 0);
    ( USERCLK *> MAXISRCTKEEP[6]) = (0, 0);
    ( USERCLK *> MAXISRCTKEEP[7]) = (0, 0);
    ( USERCLK *> MAXISRCTLAST) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[0]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[10]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[11]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[12]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[13]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[14]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[15]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[16]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[17]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[18]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[19]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[1]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[20]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[21]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[22]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[23]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[24]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[25]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[26]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[27]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[28]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[29]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[2]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[30]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[31]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[32]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[33]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[34]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[35]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[36]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[37]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[38]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[39]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[3]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[40]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[41]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[42]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[43]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[44]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[45]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[46]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[47]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[48]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[49]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[4]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[50]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[51]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[52]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[53]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[54]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[55]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[56]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[57]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[58]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[59]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[5]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[60]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[61]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[62]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[63]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[64]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[65]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[66]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[67]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[68]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[69]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[6]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[70]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[71]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[72]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[73]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[74]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[7]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[8]) = (0, 0);
    ( USERCLK *> MAXISRCTUSER[9]) = (0, 0);
    ( USERCLK *> MAXISRCTVALID) = (0, 0);
    ( USERCLK *> PCIECQNPREQCOUNT[0]) = (0, 0);
    ( USERCLK *> PCIECQNPREQCOUNT[1]) = (0, 0);
    ( USERCLK *> PCIECQNPREQCOUNT[2]) = (0, 0);
    ( USERCLK *> PCIECQNPREQCOUNT[3]) = (0, 0);
    ( USERCLK *> PCIECQNPREQCOUNT[4]) = (0, 0);
    ( USERCLK *> PCIECQNPREQCOUNT[5]) = (0, 0);
    ( USERCLK *> PCIERQSEQNUMVLD) = (0, 0);
    ( USERCLK *> PCIERQSEQNUM[0]) = (0, 0);
    ( USERCLK *> PCIERQSEQNUM[1]) = (0, 0);
    ( USERCLK *> PCIERQSEQNUM[2]) = (0, 0);
    ( USERCLK *> PCIERQSEQNUM[3]) = (0, 0);
    ( USERCLK *> PCIERQTAGAV[0]) = (0, 0);
    ( USERCLK *> PCIERQTAGAV[1]) = (0, 0);
    ( USERCLK *> PCIERQTAGVLD) = (0, 0);
    ( USERCLK *> PCIERQTAG[0]) = (0, 0);
    ( USERCLK *> PCIERQTAG[1]) = (0, 0);
    ( USERCLK *> PCIERQTAG[2]) = (0, 0);
    ( USERCLK *> PCIERQTAG[3]) = (0, 0);
    ( USERCLK *> PCIERQTAG[4]) = (0, 0);
    ( USERCLK *> PCIERQTAG[5]) = (0, 0);
    ( USERCLK *> PCIETFCNPDAV[0]) = (0, 0);
    ( USERCLK *> PCIETFCNPDAV[1]) = (0, 0);
    ( USERCLK *> PCIETFCNPHAV[0]) = (0, 0);
    ( USERCLK *> PCIETFCNPHAV[1]) = (0, 0);
    ( USERCLK *> SAXISCCTREADY[0]) = (0, 0);
    ( USERCLK *> SAXISCCTREADY[1]) = (0, 0);
    ( USERCLK *> SAXISCCTREADY[2]) = (0, 0);
    ( USERCLK *> SAXISCCTREADY[3]) = (0, 0);
    ( USERCLK *> SAXISRQTREADY[0]) = (0, 0);
    ( USERCLK *> SAXISRQTREADY[1]) = (0, 0);
    ( USERCLK *> SAXISRQTREADY[2]) = (0, 0);
    ( USERCLK *> SAXISRQTREADY[3]) = (0, 0);

    specparam PATHPULSE$ = 0;
  endspecify
endmodule

`endcelldefine
